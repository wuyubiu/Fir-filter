// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : FirSubblock



module FirSubblock (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload,
  output              io_FirOut_valid,
  input               io_FirOut_ready,
  output     [19:0]   io_FirOut_payload,
  input               clk,
  input               reset
);
  wire                multiply_io_input_ready;
  wire                multiply_io_multiplyResult_valid;
  wire       [19:0]   multiply_io_multiplyResult_payload_0;
  wire       [19:0]   multiply_io_multiplyResult_payload_1;
  wire       [19:0]   multiply_io_multiplyResult_payload_2;
  wire       [19:0]   multiply_io_multiplyResult_payload_3;
  wire       [19:0]   multiply_io_multiplyResult_payload_4;
  wire       [19:0]   multiply_io_multiplyResult_payload_5;
  wire       [19:0]   multiply_io_multiplyResult_payload_6;
  wire       [19:0]   multiply_io_multiplyResult_payload_7;
  wire       [19:0]   multiply_io_multiplyResult_payload_8;
  wire       [19:0]   multiply_io_multiplyResult_payload_9;
  wire       [19:0]   multiply_io_multiplyResult_payload_10;
  wire       [19:0]   multiply_io_multiplyResult_payload_11;
  wire       [19:0]   multiply_io_multiplyResult_payload_12;
  wire       [19:0]   multiply_io_multiplyResult_payload_13;
  wire       [19:0]   multiply_io_multiplyResult_payload_14;
  wire       [19:0]   multiply_io_multiplyResult_payload_15;
  wire       [19:0]   multiply_io_multiplyResult_payload_16;
  wire       [19:0]   multiply_io_multiplyResult_payload_17;
  wire       [19:0]   multiply_io_multiplyResult_payload_18;
  wire       [19:0]   multiply_io_multiplyResult_payload_19;
  wire       [19:0]   multiply_io_multiplyResult_payload_20;
  wire       [19:0]   multiply_io_multiplyResult_payload_21;
  wire       [19:0]   multiply_io_multiplyResult_payload_22;
  wire       [19:0]   multiply_io_multiplyResult_payload_23;
  wire       [19:0]   multiply_io_multiplyResult_payload_24;
  wire       [19:0]   multiply_io_multiplyResult_payload_25;
  wire       [19:0]   multiply_io_multiplyResult_payload_26;
  wire       [19:0]   multiply_io_multiplyResult_payload_27;
  wire       [19:0]   multiply_io_multiplyResult_payload_28;
  wire       [19:0]   multiply_io_multiplyResult_payload_29;
  wire       [19:0]   multiply_io_multiplyResult_payload_30;
  wire       [19:0]   _zz_io_FirOut_payload;
  wire       [19:0]   _zz_io_FirOut_payload_1;
  wire       [19:0]   _zz_io_FirOut_payload_2;
  wire       [19:0]   _zz_io_FirOut_payload_3;
  wire       [19:0]   _zz_io_FirOut_payload_4;
  wire       [19:0]   _zz_io_FirOut_payload_5;
  wire       [19:0]   _zz_io_FirOut_payload_6;
  wire       [19:0]   _zz_io_FirOut_payload_7;
  wire       [19:0]   _zz_io_FirOut_payload_8;
  wire       [19:0]   _zz_io_FirOut_payload_9;
  wire       [19:0]   _zz_io_FirOut_payload_10;
  wire       [19:0]   _zz_io_FirOut_payload_11;
  wire       [19:0]   _zz_io_FirOut_payload_12;
  wire       [19:0]   _zz_io_FirOut_payload_13;
  wire       [19:0]   _zz_io_FirOut_payload_14;
  wire       [19:0]   _zz_io_FirOut_payload_15;
  wire       [19:0]   _zz_io_FirOut_payload_16;
  wire       [19:0]   _zz_io_FirOut_payload_17;
  wire       [19:0]   _zz_io_FirOut_payload_18;
  wire       [19:0]   _zz_io_FirOut_payload_19;
  wire       [19:0]   _zz_io_FirOut_payload_20;
  wire       [19:0]   _zz_io_FirOut_payload_21;
  wire       [19:0]   _zz_io_FirOut_payload_22;
  wire       [19:0]   _zz_io_FirOut_payload_23;
  wire       [19:0]   _zz_io_FirOut_payload_24;
  wire       [19:0]   _zz_io_FirOut_payload_25;
  wire       [19:0]   _zz_io_FirOut_payload_26;
  wire       [19:0]   _zz_io_FirOut_payload_27;
  wire       [19:0]   _zz_io_FirOut_payload_28;

  assign _zz_io_FirOut_payload = ($signed(_zz_io_FirOut_payload_1) + $signed(_zz_io_FirOut_payload_8));
  assign _zz_io_FirOut_payload_1 = ($signed(_zz_io_FirOut_payload_2) + $signed(_zz_io_FirOut_payload_5));
  assign _zz_io_FirOut_payload_2 = ($signed(_zz_io_FirOut_payload_3) + $signed(_zz_io_FirOut_payload_4));
  assign _zz_io_FirOut_payload_3 = ($signed(multiply_io_multiplyResult_payload_0) + $signed(multiply_io_multiplyResult_payload_1));
  assign _zz_io_FirOut_payload_4 = ($signed(multiply_io_multiplyResult_payload_2) + $signed(multiply_io_multiplyResult_payload_3));
  assign _zz_io_FirOut_payload_5 = ($signed(_zz_io_FirOut_payload_6) + $signed(_zz_io_FirOut_payload_7));
  assign _zz_io_FirOut_payload_6 = ($signed(multiply_io_multiplyResult_payload_4) + $signed(multiply_io_multiplyResult_payload_5));
  assign _zz_io_FirOut_payload_7 = ($signed(multiply_io_multiplyResult_payload_6) + $signed(multiply_io_multiplyResult_payload_7));
  assign _zz_io_FirOut_payload_8 = ($signed(_zz_io_FirOut_payload_9) + $signed(_zz_io_FirOut_payload_12));
  assign _zz_io_FirOut_payload_9 = ($signed(_zz_io_FirOut_payload_10) + $signed(_zz_io_FirOut_payload_11));
  assign _zz_io_FirOut_payload_10 = ($signed(multiply_io_multiplyResult_payload_8) + $signed(multiply_io_multiplyResult_payload_9));
  assign _zz_io_FirOut_payload_11 = ($signed(multiply_io_multiplyResult_payload_10) + $signed(multiply_io_multiplyResult_payload_11));
  assign _zz_io_FirOut_payload_12 = ($signed(_zz_io_FirOut_payload_13) + $signed(_zz_io_FirOut_payload_14));
  assign _zz_io_FirOut_payload_13 = ($signed(multiply_io_multiplyResult_payload_12) + $signed(multiply_io_multiplyResult_payload_13));
  assign _zz_io_FirOut_payload_14 = ($signed(multiply_io_multiplyResult_payload_14) + $signed(multiply_io_multiplyResult_payload_15));
  assign _zz_io_FirOut_payload_15 = ($signed(_zz_io_FirOut_payload_16) + $signed(_zz_io_FirOut_payload_23));
  assign _zz_io_FirOut_payload_16 = ($signed(_zz_io_FirOut_payload_17) + $signed(_zz_io_FirOut_payload_20));
  assign _zz_io_FirOut_payload_17 = ($signed(_zz_io_FirOut_payload_18) + $signed(_zz_io_FirOut_payload_19));
  assign _zz_io_FirOut_payload_18 = ($signed(multiply_io_multiplyResult_payload_16) + $signed(multiply_io_multiplyResult_payload_17));
  assign _zz_io_FirOut_payload_19 = ($signed(multiply_io_multiplyResult_payload_18) + $signed(multiply_io_multiplyResult_payload_19));
  assign _zz_io_FirOut_payload_20 = ($signed(_zz_io_FirOut_payload_21) + $signed(_zz_io_FirOut_payload_22));
  assign _zz_io_FirOut_payload_21 = ($signed(multiply_io_multiplyResult_payload_20) + $signed(multiply_io_multiplyResult_payload_21));
  assign _zz_io_FirOut_payload_22 = ($signed(multiply_io_multiplyResult_payload_22) + $signed(multiply_io_multiplyResult_payload_23));
  assign _zz_io_FirOut_payload_23 = ($signed(_zz_io_FirOut_payload_24) + $signed(_zz_io_FirOut_payload_27));
  assign _zz_io_FirOut_payload_24 = ($signed(_zz_io_FirOut_payload_25) + $signed(_zz_io_FirOut_payload_26));
  assign _zz_io_FirOut_payload_25 = ($signed(multiply_io_multiplyResult_payload_24) + $signed(multiply_io_multiplyResult_payload_25));
  assign _zz_io_FirOut_payload_26 = ($signed(multiply_io_multiplyResult_payload_26) + $signed(multiply_io_multiplyResult_payload_27));
  assign _zz_io_FirOut_payload_27 = ($signed(_zz_io_FirOut_payload_28) + $signed(multiply_io_multiplyResult_payload_30));
  assign _zz_io_FirOut_payload_28 = ($signed(multiply_io_multiplyResult_payload_28) + $signed(multiply_io_multiplyResult_payload_29));
  MultiplyStream multiply (
    .io_input_valid                  (io_input_valid                         ), //i
    .io_input_ready                  (multiply_io_input_ready                ), //o
    .io_input_payload                (io_input_payload                       ), //i
    .io_multiplyResult_valid         (multiply_io_multiplyResult_valid       ), //o
    .io_multiplyResult_ready         (io_FirOut_ready                        ), //i
    .io_multiplyResult_payload_0     (multiply_io_multiplyResult_payload_0   ), //o
    .io_multiplyResult_payload_1     (multiply_io_multiplyResult_payload_1   ), //o
    .io_multiplyResult_payload_2     (multiply_io_multiplyResult_payload_2   ), //o
    .io_multiplyResult_payload_3     (multiply_io_multiplyResult_payload_3   ), //o
    .io_multiplyResult_payload_4     (multiply_io_multiplyResult_payload_4   ), //o
    .io_multiplyResult_payload_5     (multiply_io_multiplyResult_payload_5   ), //o
    .io_multiplyResult_payload_6     (multiply_io_multiplyResult_payload_6   ), //o
    .io_multiplyResult_payload_7     (multiply_io_multiplyResult_payload_7   ), //o
    .io_multiplyResult_payload_8     (multiply_io_multiplyResult_payload_8   ), //o
    .io_multiplyResult_payload_9     (multiply_io_multiplyResult_payload_9   ), //o
    .io_multiplyResult_payload_10    (multiply_io_multiplyResult_payload_10  ), //o
    .io_multiplyResult_payload_11    (multiply_io_multiplyResult_payload_11  ), //o
    .io_multiplyResult_payload_12    (multiply_io_multiplyResult_payload_12  ), //o
    .io_multiplyResult_payload_13    (multiply_io_multiplyResult_payload_13  ), //o
    .io_multiplyResult_payload_14    (multiply_io_multiplyResult_payload_14  ), //o
    .io_multiplyResult_payload_15    (multiply_io_multiplyResult_payload_15  ), //o
    .io_multiplyResult_payload_16    (multiply_io_multiplyResult_payload_16  ), //o
    .io_multiplyResult_payload_17    (multiply_io_multiplyResult_payload_17  ), //o
    .io_multiplyResult_payload_18    (multiply_io_multiplyResult_payload_18  ), //o
    .io_multiplyResult_payload_19    (multiply_io_multiplyResult_payload_19  ), //o
    .io_multiplyResult_payload_20    (multiply_io_multiplyResult_payload_20  ), //o
    .io_multiplyResult_payload_21    (multiply_io_multiplyResult_payload_21  ), //o
    .io_multiplyResult_payload_22    (multiply_io_multiplyResult_payload_22  ), //o
    .io_multiplyResult_payload_23    (multiply_io_multiplyResult_payload_23  ), //o
    .io_multiplyResult_payload_24    (multiply_io_multiplyResult_payload_24  ), //o
    .io_multiplyResult_payload_25    (multiply_io_multiplyResult_payload_25  ), //o
    .io_multiplyResult_payload_26    (multiply_io_multiplyResult_payload_26  ), //o
    .io_multiplyResult_payload_27    (multiply_io_multiplyResult_payload_27  ), //o
    .io_multiplyResult_payload_28    (multiply_io_multiplyResult_payload_28  ), //o
    .io_multiplyResult_payload_29    (multiply_io_multiplyResult_payload_29  ), //o
    .io_multiplyResult_payload_30    (multiply_io_multiplyResult_payload_30  ), //o
    .clk                             (clk                                    ), //i
    .reset                           (reset                                  )  //i
  );
  assign io_input_ready = multiply_io_input_ready;
  assign io_FirOut_valid = multiply_io_multiplyResult_valid;
  assign io_FirOut_payload = ($signed(_zz_io_FirOut_payload) + $signed(_zz_io_FirOut_payload_15));

endmodule

module MultiplyStream (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload,
  output              io_multiplyResult_valid,
  input               io_multiplyResult_ready,
  output     [19:0]   io_multiplyResult_payload_0,
  output     [19:0]   io_multiplyResult_payload_1,
  output     [19:0]   io_multiplyResult_payload_2,
  output     [19:0]   io_multiplyResult_payload_3,
  output     [19:0]   io_multiplyResult_payload_4,
  output     [19:0]   io_multiplyResult_payload_5,
  output     [19:0]   io_multiplyResult_payload_6,
  output     [19:0]   io_multiplyResult_payload_7,
  output     [19:0]   io_multiplyResult_payload_8,
  output     [19:0]   io_multiplyResult_payload_9,
  output     [19:0]   io_multiplyResult_payload_10,
  output     [19:0]   io_multiplyResult_payload_11,
  output     [19:0]   io_multiplyResult_payload_12,
  output     [19:0]   io_multiplyResult_payload_13,
  output     [19:0]   io_multiplyResult_payload_14,
  output     [19:0]   io_multiplyResult_payload_15,
  output     [19:0]   io_multiplyResult_payload_16,
  output     [19:0]   io_multiplyResult_payload_17,
  output     [19:0]   io_multiplyResult_payload_18,
  output     [19:0]   io_multiplyResult_payload_19,
  output     [19:0]   io_multiplyResult_payload_20,
  output     [19:0]   io_multiplyResult_payload_21,
  output     [19:0]   io_multiplyResult_payload_22,
  output     [19:0]   io_multiplyResult_payload_23,
  output     [19:0]   io_multiplyResult_payload_24,
  output     [19:0]   io_multiplyResult_payload_25,
  output     [19:0]   io_multiplyResult_payload_26,
  output     [19:0]   io_multiplyResult_payload_27,
  output     [19:0]   io_multiplyResult_payload_28,
  output     [19:0]   io_multiplyResult_payload_29,
  output     [19:0]   io_multiplyResult_payload_30,
  input               clk,
  input               reset
);
  reg                 signalInput_0_fork_io_outputs_0_ready;
  reg                 signalInput_1_fork_io_outputs_0_ready;
  reg                 signalInput_2_fork_io_outputs_0_ready;
  reg                 signalInput_3_fork_io_outputs_0_ready;
  reg                 signalInput_4_fork_io_outputs_0_ready;
  reg                 signalInput_5_fork_io_outputs_0_ready;
  reg                 signalInput_6_fork_io_outputs_0_ready;
  reg                 signalInput_7_fork_io_outputs_0_ready;
  reg                 signalInput_8_fork_io_outputs_0_ready;
  reg                 signalInput_9_fork_io_outputs_0_ready;
  reg                 signalInput_10_fork_io_outputs_0_ready;
  reg                 signalInput_11_fork_io_outputs_0_ready;
  reg                 signalInput_12_fork_io_outputs_0_ready;
  reg                 signalInput_13_fork_io_outputs_0_ready;
  reg                 signalInput_14_fork_io_outputs_0_ready;
  reg                 signalInput_15_fork_io_outputs_0_ready;
  reg                 signalInput_16_fork_io_outputs_0_ready;
  reg                 signalInput_17_fork_io_outputs_0_ready;
  reg                 signalInput_18_fork_io_outputs_0_ready;
  reg                 signalInput_19_fork_io_outputs_0_ready;
  reg                 signalInput_20_fork_io_outputs_0_ready;
  reg                 signalInput_21_fork_io_outputs_0_ready;
  reg                 signalInput_22_fork_io_outputs_0_ready;
  reg                 signalInput_23_fork_io_outputs_0_ready;
  reg                 signalInput_24_fork_io_outputs_0_ready;
  reg                 signalInput_25_fork_io_outputs_0_ready;
  reg                 signalInput_26_fork_io_outputs_0_ready;
  reg                 signalInput_27_fork_io_outputs_0_ready;
  reg                 signalInput_28_fork_io_outputs_0_ready;
  reg                 signalInput_29_fork_io_outputs_0_ready;
  reg                 signalInput_30_fork_io_outputs_0_ready;
  wire                signalInput_0_fork_io_input_ready;
  wire                signalInput_0_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_0_fork_io_outputs_0_payload;
  wire                signalInput_0_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_0_fork_io_outputs_1_payload;
  wire                signalInput_1_fork_io_input_ready;
  wire                signalInput_1_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_1_fork_io_outputs_0_payload;
  wire                signalInput_1_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_1_fork_io_outputs_1_payload;
  wire                signalInput_2_fork_io_input_ready;
  wire                signalInput_2_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_2_fork_io_outputs_0_payload;
  wire                signalInput_2_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_2_fork_io_outputs_1_payload;
  wire                signalInput_3_fork_io_input_ready;
  wire                signalInput_3_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_3_fork_io_outputs_0_payload;
  wire                signalInput_3_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_3_fork_io_outputs_1_payload;
  wire                signalInput_4_fork_io_input_ready;
  wire                signalInput_4_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_4_fork_io_outputs_0_payload;
  wire                signalInput_4_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_4_fork_io_outputs_1_payload;
  wire                signalInput_5_fork_io_input_ready;
  wire                signalInput_5_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_5_fork_io_outputs_0_payload;
  wire                signalInput_5_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_5_fork_io_outputs_1_payload;
  wire                signalInput_6_fork_io_input_ready;
  wire                signalInput_6_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_6_fork_io_outputs_0_payload;
  wire                signalInput_6_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_6_fork_io_outputs_1_payload;
  wire                signalInput_7_fork_io_input_ready;
  wire                signalInput_7_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_7_fork_io_outputs_0_payload;
  wire                signalInput_7_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_7_fork_io_outputs_1_payload;
  wire                signalInput_8_fork_io_input_ready;
  wire                signalInput_8_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_8_fork_io_outputs_0_payload;
  wire                signalInput_8_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_8_fork_io_outputs_1_payload;
  wire                signalInput_9_fork_io_input_ready;
  wire                signalInput_9_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_9_fork_io_outputs_0_payload;
  wire                signalInput_9_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_9_fork_io_outputs_1_payload;
  wire                signalInput_10_fork_io_input_ready;
  wire                signalInput_10_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_10_fork_io_outputs_0_payload;
  wire                signalInput_10_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_10_fork_io_outputs_1_payload;
  wire                signalInput_11_fork_io_input_ready;
  wire                signalInput_11_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_11_fork_io_outputs_0_payload;
  wire                signalInput_11_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_11_fork_io_outputs_1_payload;
  wire                signalInput_12_fork_io_input_ready;
  wire                signalInput_12_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_12_fork_io_outputs_0_payload;
  wire                signalInput_12_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_12_fork_io_outputs_1_payload;
  wire                signalInput_13_fork_io_input_ready;
  wire                signalInput_13_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_13_fork_io_outputs_0_payload;
  wire                signalInput_13_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_13_fork_io_outputs_1_payload;
  wire                signalInput_14_fork_io_input_ready;
  wire                signalInput_14_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_14_fork_io_outputs_0_payload;
  wire                signalInput_14_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_14_fork_io_outputs_1_payload;
  wire                signalInput_15_fork_io_input_ready;
  wire                signalInput_15_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_15_fork_io_outputs_0_payload;
  wire                signalInput_15_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_15_fork_io_outputs_1_payload;
  wire                signalInput_16_fork_io_input_ready;
  wire                signalInput_16_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_16_fork_io_outputs_0_payload;
  wire                signalInput_16_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_16_fork_io_outputs_1_payload;
  wire                signalInput_17_fork_io_input_ready;
  wire                signalInput_17_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_17_fork_io_outputs_0_payload;
  wire                signalInput_17_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_17_fork_io_outputs_1_payload;
  wire                signalInput_18_fork_io_input_ready;
  wire                signalInput_18_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_18_fork_io_outputs_0_payload;
  wire                signalInput_18_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_18_fork_io_outputs_1_payload;
  wire                signalInput_19_fork_io_input_ready;
  wire                signalInput_19_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_19_fork_io_outputs_0_payload;
  wire                signalInput_19_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_19_fork_io_outputs_1_payload;
  wire                signalInput_20_fork_io_input_ready;
  wire                signalInput_20_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_20_fork_io_outputs_0_payload;
  wire                signalInput_20_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_20_fork_io_outputs_1_payload;
  wire                signalInput_21_fork_io_input_ready;
  wire                signalInput_21_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_21_fork_io_outputs_0_payload;
  wire                signalInput_21_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_21_fork_io_outputs_1_payload;
  wire                signalInput_22_fork_io_input_ready;
  wire                signalInput_22_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_22_fork_io_outputs_0_payload;
  wire                signalInput_22_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_22_fork_io_outputs_1_payload;
  wire                signalInput_23_fork_io_input_ready;
  wire                signalInput_23_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_23_fork_io_outputs_0_payload;
  wire                signalInput_23_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_23_fork_io_outputs_1_payload;
  wire                signalInput_24_fork_io_input_ready;
  wire                signalInput_24_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_24_fork_io_outputs_0_payload;
  wire                signalInput_24_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_24_fork_io_outputs_1_payload;
  wire                signalInput_25_fork_io_input_ready;
  wire                signalInput_25_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_25_fork_io_outputs_0_payload;
  wire                signalInput_25_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_25_fork_io_outputs_1_payload;
  wire                signalInput_26_fork_io_input_ready;
  wire                signalInput_26_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_26_fork_io_outputs_0_payload;
  wire                signalInput_26_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_26_fork_io_outputs_1_payload;
  wire                signalInput_27_fork_io_input_ready;
  wire                signalInput_27_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_27_fork_io_outputs_0_payload;
  wire                signalInput_27_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_27_fork_io_outputs_1_payload;
  wire                signalInput_28_fork_io_input_ready;
  wire                signalInput_28_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_28_fork_io_outputs_0_payload;
  wire                signalInput_28_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_28_fork_io_outputs_1_payload;
  wire                signalInput_29_fork_io_input_ready;
  wire                signalInput_29_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_29_fork_io_outputs_0_payload;
  wire                signalInput_29_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_29_fork_io_outputs_1_payload;
  wire                signalInput_30_fork_io_input_ready;
  wire                signalInput_30_fork_io_outputs_0_valid;
  wire       [7:0]    signalInput_30_fork_io_outputs_0_payload;
  wire                signalInput_30_fork_io_outputs_1_valid;
  wire       [7:0]    signalInput_30_fork_io_outputs_1_payload;
  wire       [16:0]   _zz_signalInput_0_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_0_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_1_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_1_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_2_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_2_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_3_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_3_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_4_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_4_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_5_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_5_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_6_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_6_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_7_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_7_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_8_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_8_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_9_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_9_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_10_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_10_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_11_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_11_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_12_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_12_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_13_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_13_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_14_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_14_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_15_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_15_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_16_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_16_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_17_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_17_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_18_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_18_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_19_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_19_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_20_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_20_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_21_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_21_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_22_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_22_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_23_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_23_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_24_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_24_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_25_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_25_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_26_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_26_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_27_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_27_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_28_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_28_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_29_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_29_fork_io_outputs_1_translated_payload_1;
  wire       [16:0]   _zz_signalInput_30_fork_io_outputs_1_translated_payload;
  wire       [8:0]    _zz_signalInput_30_fork_io_outputs_1_translated_payload_1;
  wire                _zz_io_multiplyResult_valid;
  wire                signalInput_0_valid;
  wire                signalInput_0_ready;
  wire       [7:0]    signalInput_0_payload;
  wire                signalInput_1_valid;
  wire                signalInput_1_ready;
  wire       [7:0]    signalInput_1_payload;
  wire                signalInput_2_valid;
  wire                signalInput_2_ready;
  wire       [7:0]    signalInput_2_payload;
  wire                signalInput_3_valid;
  wire                signalInput_3_ready;
  wire       [7:0]    signalInput_3_payload;
  wire                signalInput_4_valid;
  wire                signalInput_4_ready;
  wire       [7:0]    signalInput_4_payload;
  wire                signalInput_5_valid;
  wire                signalInput_5_ready;
  wire       [7:0]    signalInput_5_payload;
  wire                signalInput_6_valid;
  wire                signalInput_6_ready;
  wire       [7:0]    signalInput_6_payload;
  wire                signalInput_7_valid;
  wire                signalInput_7_ready;
  wire       [7:0]    signalInput_7_payload;
  wire                signalInput_8_valid;
  wire                signalInput_8_ready;
  wire       [7:0]    signalInput_8_payload;
  wire                signalInput_9_valid;
  wire                signalInput_9_ready;
  wire       [7:0]    signalInput_9_payload;
  wire                signalInput_10_valid;
  wire                signalInput_10_ready;
  wire       [7:0]    signalInput_10_payload;
  wire                signalInput_11_valid;
  wire                signalInput_11_ready;
  wire       [7:0]    signalInput_11_payload;
  wire                signalInput_12_valid;
  wire                signalInput_12_ready;
  wire       [7:0]    signalInput_12_payload;
  wire                signalInput_13_valid;
  wire                signalInput_13_ready;
  wire       [7:0]    signalInput_13_payload;
  wire                signalInput_14_valid;
  wire                signalInput_14_ready;
  wire       [7:0]    signalInput_14_payload;
  wire                signalInput_15_valid;
  wire                signalInput_15_ready;
  wire       [7:0]    signalInput_15_payload;
  wire                signalInput_16_valid;
  wire                signalInput_16_ready;
  wire       [7:0]    signalInput_16_payload;
  wire                signalInput_17_valid;
  wire                signalInput_17_ready;
  wire       [7:0]    signalInput_17_payload;
  wire                signalInput_18_valid;
  wire                signalInput_18_ready;
  wire       [7:0]    signalInput_18_payload;
  wire                signalInput_19_valid;
  wire                signalInput_19_ready;
  wire       [7:0]    signalInput_19_payload;
  wire                signalInput_20_valid;
  wire                signalInput_20_ready;
  wire       [7:0]    signalInput_20_payload;
  wire                signalInput_21_valid;
  wire                signalInput_21_ready;
  wire       [7:0]    signalInput_21_payload;
  wire                signalInput_22_valid;
  wire                signalInput_22_ready;
  wire       [7:0]    signalInput_22_payload;
  wire                signalInput_23_valid;
  wire                signalInput_23_ready;
  wire       [7:0]    signalInput_23_payload;
  wire                signalInput_24_valid;
  wire                signalInput_24_ready;
  wire       [7:0]    signalInput_24_payload;
  wire                signalInput_25_valid;
  wire                signalInput_25_ready;
  wire       [7:0]    signalInput_25_payload;
  wire                signalInput_26_valid;
  wire                signalInput_26_ready;
  wire       [7:0]    signalInput_26_payload;
  wire                signalInput_27_valid;
  wire                signalInput_27_ready;
  wire       [7:0]    signalInput_27_payload;
  wire                signalInput_28_valid;
  wire                signalInput_28_ready;
  wire       [7:0]    signalInput_28_payload;
  wire                signalInput_29_valid;
  wire                signalInput_29_ready;
  wire       [7:0]    signalInput_29_payload;
  wire                signalInput_30_valid;
  wire                signalInput_30_ready;
  wire       [7:0]    signalInput_30_payload;
  wire                mulOut_0_valid;
  wire                mulOut_0_ready;
  wire       [19:0]   mulOut_0_payload;
  wire                signalInput_0_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_0_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_0_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_0_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_0_fork_io_outputs_0_rData;
  wire                when_Stream_l342;
  wire                signalInput_0_fork_io_outputs_1_translated_valid;
  wire                signalInput_0_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_0_fork_io_outputs_1_translated_payload;
  wire                mulOut_1_valid;
  wire                mulOut_1_ready;
  wire       [19:0]   mulOut_1_payload;
  wire                signalInput_1_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_1_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_1_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_1_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_1_fork_io_outputs_0_rData;
  wire                when_Stream_l342_1;
  wire                signalInput_1_fork_io_outputs_1_translated_valid;
  wire                signalInput_1_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_1_fork_io_outputs_1_translated_payload;
  wire                mulOut_2_valid;
  wire                mulOut_2_ready;
  wire       [19:0]   mulOut_2_payload;
  wire                signalInput_2_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_2_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_2_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_2_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_2_fork_io_outputs_0_rData;
  wire                when_Stream_l342_2;
  wire                signalInput_2_fork_io_outputs_1_translated_valid;
  wire                signalInput_2_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_2_fork_io_outputs_1_translated_payload;
  wire                mulOut_3_valid;
  wire                mulOut_3_ready;
  wire       [19:0]   mulOut_3_payload;
  wire                signalInput_3_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_3_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_3_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_3_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_3_fork_io_outputs_0_rData;
  wire                when_Stream_l342_3;
  wire                signalInput_3_fork_io_outputs_1_translated_valid;
  wire                signalInput_3_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_3_fork_io_outputs_1_translated_payload;
  wire                mulOut_4_valid;
  wire                mulOut_4_ready;
  wire       [19:0]   mulOut_4_payload;
  wire                signalInput_4_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_4_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_4_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_4_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_4_fork_io_outputs_0_rData;
  wire                when_Stream_l342_4;
  wire                signalInput_4_fork_io_outputs_1_translated_valid;
  wire                signalInput_4_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_4_fork_io_outputs_1_translated_payload;
  wire                mulOut_5_valid;
  wire                mulOut_5_ready;
  wire       [19:0]   mulOut_5_payload;
  wire                signalInput_5_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_5_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_5_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_5_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_5_fork_io_outputs_0_rData;
  wire                when_Stream_l342_5;
  wire                signalInput_5_fork_io_outputs_1_translated_valid;
  wire                signalInput_5_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_5_fork_io_outputs_1_translated_payload;
  wire                mulOut_6_valid;
  wire                mulOut_6_ready;
  wire       [19:0]   mulOut_6_payload;
  wire                signalInput_6_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_6_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_6_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_6_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_6_fork_io_outputs_0_rData;
  wire                when_Stream_l342_6;
  wire                signalInput_6_fork_io_outputs_1_translated_valid;
  wire                signalInput_6_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_6_fork_io_outputs_1_translated_payload;
  wire                mulOut_7_valid;
  wire                mulOut_7_ready;
  wire       [19:0]   mulOut_7_payload;
  wire                signalInput_7_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_7_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_7_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_7_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_7_fork_io_outputs_0_rData;
  wire                when_Stream_l342_7;
  wire                signalInput_7_fork_io_outputs_1_translated_valid;
  wire                signalInput_7_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_7_fork_io_outputs_1_translated_payload;
  wire                mulOut_8_valid;
  wire                mulOut_8_ready;
  wire       [19:0]   mulOut_8_payload;
  wire                signalInput_8_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_8_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_8_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_8_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_8_fork_io_outputs_0_rData;
  wire                when_Stream_l342_8;
  wire                signalInput_8_fork_io_outputs_1_translated_valid;
  wire                signalInput_8_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_8_fork_io_outputs_1_translated_payload;
  wire                mulOut_9_valid;
  wire                mulOut_9_ready;
  wire       [19:0]   mulOut_9_payload;
  wire                signalInput_9_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_9_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_9_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_9_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_9_fork_io_outputs_0_rData;
  wire                when_Stream_l342_9;
  wire                signalInput_9_fork_io_outputs_1_translated_valid;
  wire                signalInput_9_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_9_fork_io_outputs_1_translated_payload;
  wire                mulOut_10_valid;
  wire                mulOut_10_ready;
  wire       [19:0]   mulOut_10_payload;
  wire                signalInput_10_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_10_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_10_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_10_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_10_fork_io_outputs_0_rData;
  wire                when_Stream_l342_10;
  wire                signalInput_10_fork_io_outputs_1_translated_valid;
  wire                signalInput_10_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_10_fork_io_outputs_1_translated_payload;
  wire                mulOut_11_valid;
  wire                mulOut_11_ready;
  wire       [19:0]   mulOut_11_payload;
  wire                signalInput_11_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_11_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_11_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_11_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_11_fork_io_outputs_0_rData;
  wire                when_Stream_l342_11;
  wire                signalInput_11_fork_io_outputs_1_translated_valid;
  wire                signalInput_11_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_11_fork_io_outputs_1_translated_payload;
  wire                mulOut_12_valid;
  wire                mulOut_12_ready;
  wire       [19:0]   mulOut_12_payload;
  wire                signalInput_12_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_12_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_12_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_12_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_12_fork_io_outputs_0_rData;
  wire                when_Stream_l342_12;
  wire                signalInput_12_fork_io_outputs_1_translated_valid;
  wire                signalInput_12_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_12_fork_io_outputs_1_translated_payload;
  wire                mulOut_13_valid;
  wire                mulOut_13_ready;
  wire       [19:0]   mulOut_13_payload;
  wire                signalInput_13_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_13_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_13_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_13_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_13_fork_io_outputs_0_rData;
  wire                when_Stream_l342_13;
  wire                signalInput_13_fork_io_outputs_1_translated_valid;
  wire                signalInput_13_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_13_fork_io_outputs_1_translated_payload;
  wire                mulOut_14_valid;
  wire                mulOut_14_ready;
  wire       [19:0]   mulOut_14_payload;
  wire                signalInput_14_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_14_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_14_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_14_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_14_fork_io_outputs_0_rData;
  wire                when_Stream_l342_14;
  wire                signalInput_14_fork_io_outputs_1_translated_valid;
  wire                signalInput_14_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_14_fork_io_outputs_1_translated_payload;
  wire                mulOut_15_valid;
  wire                mulOut_15_ready;
  wire       [19:0]   mulOut_15_payload;
  wire                signalInput_15_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_15_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_15_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_15_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_15_fork_io_outputs_0_rData;
  wire                when_Stream_l342_15;
  wire                signalInput_15_fork_io_outputs_1_translated_valid;
  wire                signalInput_15_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_15_fork_io_outputs_1_translated_payload;
  wire                mulOut_16_valid;
  wire                mulOut_16_ready;
  wire       [19:0]   mulOut_16_payload;
  wire                signalInput_16_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_16_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_16_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_16_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_16_fork_io_outputs_0_rData;
  wire                when_Stream_l342_16;
  wire                signalInput_16_fork_io_outputs_1_translated_valid;
  wire                signalInput_16_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_16_fork_io_outputs_1_translated_payload;
  wire                mulOut_17_valid;
  wire                mulOut_17_ready;
  wire       [19:0]   mulOut_17_payload;
  wire                signalInput_17_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_17_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_17_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_17_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_17_fork_io_outputs_0_rData;
  wire                when_Stream_l342_17;
  wire                signalInput_17_fork_io_outputs_1_translated_valid;
  wire                signalInput_17_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_17_fork_io_outputs_1_translated_payload;
  wire                mulOut_18_valid;
  wire                mulOut_18_ready;
  wire       [19:0]   mulOut_18_payload;
  wire                signalInput_18_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_18_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_18_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_18_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_18_fork_io_outputs_0_rData;
  wire                when_Stream_l342_18;
  wire                signalInput_18_fork_io_outputs_1_translated_valid;
  wire                signalInput_18_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_18_fork_io_outputs_1_translated_payload;
  wire                mulOut_19_valid;
  wire                mulOut_19_ready;
  wire       [19:0]   mulOut_19_payload;
  wire                signalInput_19_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_19_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_19_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_19_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_19_fork_io_outputs_0_rData;
  wire                when_Stream_l342_19;
  wire                signalInput_19_fork_io_outputs_1_translated_valid;
  wire                signalInput_19_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_19_fork_io_outputs_1_translated_payload;
  wire                mulOut_20_valid;
  wire                mulOut_20_ready;
  wire       [19:0]   mulOut_20_payload;
  wire                signalInput_20_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_20_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_20_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_20_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_20_fork_io_outputs_0_rData;
  wire                when_Stream_l342_20;
  wire                signalInput_20_fork_io_outputs_1_translated_valid;
  wire                signalInput_20_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_20_fork_io_outputs_1_translated_payload;
  wire                mulOut_21_valid;
  wire                mulOut_21_ready;
  wire       [19:0]   mulOut_21_payload;
  wire                signalInput_21_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_21_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_21_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_21_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_21_fork_io_outputs_0_rData;
  wire                when_Stream_l342_21;
  wire                signalInput_21_fork_io_outputs_1_translated_valid;
  wire                signalInput_21_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_21_fork_io_outputs_1_translated_payload;
  wire                mulOut_22_valid;
  wire                mulOut_22_ready;
  wire       [19:0]   mulOut_22_payload;
  wire                signalInput_22_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_22_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_22_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_22_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_22_fork_io_outputs_0_rData;
  wire                when_Stream_l342_22;
  wire                signalInput_22_fork_io_outputs_1_translated_valid;
  wire                signalInput_22_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_22_fork_io_outputs_1_translated_payload;
  wire                mulOut_23_valid;
  wire                mulOut_23_ready;
  wire       [19:0]   mulOut_23_payload;
  wire                signalInput_23_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_23_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_23_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_23_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_23_fork_io_outputs_0_rData;
  wire                when_Stream_l342_23;
  wire                signalInput_23_fork_io_outputs_1_translated_valid;
  wire                signalInput_23_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_23_fork_io_outputs_1_translated_payload;
  wire                mulOut_24_valid;
  wire                mulOut_24_ready;
  wire       [19:0]   mulOut_24_payload;
  wire                signalInput_24_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_24_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_24_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_24_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_24_fork_io_outputs_0_rData;
  wire                when_Stream_l342_24;
  wire                signalInput_24_fork_io_outputs_1_translated_valid;
  wire                signalInput_24_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_24_fork_io_outputs_1_translated_payload;
  wire                mulOut_25_valid;
  wire                mulOut_25_ready;
  wire       [19:0]   mulOut_25_payload;
  wire                signalInput_25_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_25_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_25_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_25_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_25_fork_io_outputs_0_rData;
  wire                when_Stream_l342_25;
  wire                signalInput_25_fork_io_outputs_1_translated_valid;
  wire                signalInput_25_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_25_fork_io_outputs_1_translated_payload;
  wire                mulOut_26_valid;
  wire                mulOut_26_ready;
  wire       [19:0]   mulOut_26_payload;
  wire                signalInput_26_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_26_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_26_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_26_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_26_fork_io_outputs_0_rData;
  wire                when_Stream_l342_26;
  wire                signalInput_26_fork_io_outputs_1_translated_valid;
  wire                signalInput_26_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_26_fork_io_outputs_1_translated_payload;
  wire                mulOut_27_valid;
  wire                mulOut_27_ready;
  wire       [19:0]   mulOut_27_payload;
  wire                signalInput_27_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_27_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_27_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_27_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_27_fork_io_outputs_0_rData;
  wire                when_Stream_l342_27;
  wire                signalInput_27_fork_io_outputs_1_translated_valid;
  wire                signalInput_27_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_27_fork_io_outputs_1_translated_payload;
  wire                mulOut_28_valid;
  wire                mulOut_28_ready;
  wire       [19:0]   mulOut_28_payload;
  wire                signalInput_28_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_28_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_28_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_28_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_28_fork_io_outputs_0_rData;
  wire                when_Stream_l342_28;
  wire                signalInput_28_fork_io_outputs_1_translated_valid;
  wire                signalInput_28_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_28_fork_io_outputs_1_translated_payload;
  wire                mulOut_29_valid;
  wire                mulOut_29_ready;
  wire       [19:0]   mulOut_29_payload;
  wire                signalInput_29_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_29_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_29_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_29_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_29_fork_io_outputs_0_rData;
  wire                when_Stream_l342_29;
  wire                signalInput_29_fork_io_outputs_1_translated_valid;
  wire                signalInput_29_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_29_fork_io_outputs_1_translated_payload;
  wire                mulOut_30_valid;
  wire                mulOut_30_ready;
  wire       [19:0]   mulOut_30_payload;
  wire                signalInput_30_fork_io_outputs_0_m2sPipe_valid;
  wire                signalInput_30_fork_io_outputs_0_m2sPipe_ready;
  wire       [7:0]    signalInput_30_fork_io_outputs_0_m2sPipe_payload;
  reg                 signalInput_30_fork_io_outputs_0_rValid;
  reg        [7:0]    signalInput_30_fork_io_outputs_0_rData;
  wire                when_Stream_l342_30;
  wire                signalInput_30_fork_io_outputs_1_translated_valid;
  wire                signalInput_30_fork_io_outputs_1_translated_ready;
  wire       [19:0]   signalInput_30_fork_io_outputs_1_translated_payload;

  assign _zz_signalInput_0_fork_io_outputs_1_translated_payload = ($signed(signalInput_0_fork_io_outputs_1_payload) * $signed(_zz_signalInput_0_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_0_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_1_fork_io_outputs_1_translated_payload = ($signed(signalInput_1_fork_io_outputs_1_payload) * $signed(_zz_signalInput_1_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_1_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_2_fork_io_outputs_1_translated_payload = ($signed(signalInput_2_fork_io_outputs_1_payload) * $signed(_zz_signalInput_2_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_2_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_3_fork_io_outputs_1_translated_payload = ($signed(signalInput_3_fork_io_outputs_1_payload) * $signed(_zz_signalInput_3_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_3_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_4_fork_io_outputs_1_translated_payload = ($signed(signalInput_4_fork_io_outputs_1_payload) * $signed(_zz_signalInput_4_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_4_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_5_fork_io_outputs_1_translated_payload = ($signed(signalInput_5_fork_io_outputs_1_payload) * $signed(_zz_signalInput_5_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_5_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_6_fork_io_outputs_1_translated_payload = ($signed(signalInput_6_fork_io_outputs_1_payload) * $signed(_zz_signalInput_6_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_6_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_7_fork_io_outputs_1_translated_payload = ($signed(signalInput_7_fork_io_outputs_1_payload) * $signed(_zz_signalInput_7_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_7_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_8_fork_io_outputs_1_translated_payload = ($signed(signalInput_8_fork_io_outputs_1_payload) * $signed(_zz_signalInput_8_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_8_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_9_fork_io_outputs_1_translated_payload = ($signed(signalInput_9_fork_io_outputs_1_payload) * $signed(_zz_signalInput_9_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_9_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_10_fork_io_outputs_1_translated_payload = ($signed(signalInput_10_fork_io_outputs_1_payload) * $signed(_zz_signalInput_10_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_10_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_11_fork_io_outputs_1_translated_payload = ($signed(signalInput_11_fork_io_outputs_1_payload) * $signed(_zz_signalInput_11_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_11_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_12_fork_io_outputs_1_translated_payload = ($signed(signalInput_12_fork_io_outputs_1_payload) * $signed(_zz_signalInput_12_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_12_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_13_fork_io_outputs_1_translated_payload = ($signed(signalInput_13_fork_io_outputs_1_payload) * $signed(_zz_signalInput_13_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_13_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_14_fork_io_outputs_1_translated_payload = ($signed(signalInput_14_fork_io_outputs_1_payload) * $signed(_zz_signalInput_14_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_14_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_15_fork_io_outputs_1_translated_payload = ($signed(signalInput_15_fork_io_outputs_1_payload) * $signed(_zz_signalInput_15_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_15_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_16_fork_io_outputs_1_translated_payload = ($signed(signalInput_16_fork_io_outputs_1_payload) * $signed(_zz_signalInput_16_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_16_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_17_fork_io_outputs_1_translated_payload = ($signed(signalInput_17_fork_io_outputs_1_payload) * $signed(_zz_signalInput_17_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_17_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_18_fork_io_outputs_1_translated_payload = ($signed(signalInput_18_fork_io_outputs_1_payload) * $signed(_zz_signalInput_18_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_18_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_19_fork_io_outputs_1_translated_payload = ($signed(signalInput_19_fork_io_outputs_1_payload) * $signed(_zz_signalInput_19_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_19_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_20_fork_io_outputs_1_translated_payload = ($signed(signalInput_20_fork_io_outputs_1_payload) * $signed(_zz_signalInput_20_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_20_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_21_fork_io_outputs_1_translated_payload = ($signed(signalInput_21_fork_io_outputs_1_payload) * $signed(_zz_signalInput_21_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_21_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_22_fork_io_outputs_1_translated_payload = ($signed(signalInput_22_fork_io_outputs_1_payload) * $signed(_zz_signalInput_22_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_22_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_23_fork_io_outputs_1_translated_payload = ($signed(signalInput_23_fork_io_outputs_1_payload) * $signed(_zz_signalInput_23_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_23_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_24_fork_io_outputs_1_translated_payload = ($signed(signalInput_24_fork_io_outputs_1_payload) * $signed(_zz_signalInput_24_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_24_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_25_fork_io_outputs_1_translated_payload = ($signed(signalInput_25_fork_io_outputs_1_payload) * $signed(_zz_signalInput_25_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_25_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_26_fork_io_outputs_1_translated_payload = ($signed(signalInput_26_fork_io_outputs_1_payload) * $signed(_zz_signalInput_26_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_26_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_27_fork_io_outputs_1_translated_payload = ($signed(signalInput_27_fork_io_outputs_1_payload) * $signed(_zz_signalInput_27_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_27_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_28_fork_io_outputs_1_translated_payload = ($signed(signalInput_28_fork_io_outputs_1_payload) * $signed(_zz_signalInput_28_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_28_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_29_fork_io_outputs_1_translated_payload = ($signed(signalInput_29_fork_io_outputs_1_payload) * $signed(_zz_signalInput_29_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_29_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_signalInput_30_fork_io_outputs_1_translated_payload = ($signed(signalInput_30_fork_io_outputs_1_payload) * $signed(_zz_signalInput_30_fork_io_outputs_1_translated_payload_1));
  assign _zz_signalInput_30_fork_io_outputs_1_translated_payload_1 = 9'h080;
  assign _zz_io_multiplyResult_valid = ((((((((((((((mulOut_0_valid && mulOut_1_valid) && mulOut_2_valid) && mulOut_3_valid) && mulOut_4_valid) && mulOut_5_valid) && mulOut_6_valid) && mulOut_7_valid) && mulOut_8_valid) && mulOut_9_valid) && mulOut_10_valid) && mulOut_11_valid) && mulOut_12_valid) && mulOut_13_valid) && mulOut_14_valid);
  StreamFork signalInput_0_fork (
    .io_input_valid          (signalInput_0_valid                               ), //i
    .io_input_ready          (signalInput_0_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_0_payload                             ), //i
    .io_outputs_0_valid      (signalInput_0_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_0_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_0_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_0_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_0_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_0_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_1_fork (
    .io_input_valid          (signalInput_1_valid                               ), //i
    .io_input_ready          (signalInput_1_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_1_payload                             ), //i
    .io_outputs_0_valid      (signalInput_1_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_1_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_1_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_1_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_1_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_1_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_2_fork (
    .io_input_valid          (signalInput_2_valid                               ), //i
    .io_input_ready          (signalInput_2_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_2_payload                             ), //i
    .io_outputs_0_valid      (signalInput_2_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_2_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_2_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_2_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_2_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_2_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_3_fork (
    .io_input_valid          (signalInput_3_valid                               ), //i
    .io_input_ready          (signalInput_3_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_3_payload                             ), //i
    .io_outputs_0_valid      (signalInput_3_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_3_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_3_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_3_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_3_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_3_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_4_fork (
    .io_input_valid          (signalInput_4_valid                               ), //i
    .io_input_ready          (signalInput_4_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_4_payload                             ), //i
    .io_outputs_0_valid      (signalInput_4_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_4_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_4_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_4_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_4_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_4_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_5_fork (
    .io_input_valid          (signalInput_5_valid                               ), //i
    .io_input_ready          (signalInput_5_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_5_payload                             ), //i
    .io_outputs_0_valid      (signalInput_5_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_5_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_5_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_5_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_5_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_5_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_6_fork (
    .io_input_valid          (signalInput_6_valid                               ), //i
    .io_input_ready          (signalInput_6_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_6_payload                             ), //i
    .io_outputs_0_valid      (signalInput_6_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_6_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_6_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_6_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_6_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_6_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_7_fork (
    .io_input_valid          (signalInput_7_valid                               ), //i
    .io_input_ready          (signalInput_7_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_7_payload                             ), //i
    .io_outputs_0_valid      (signalInput_7_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_7_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_7_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_7_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_7_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_7_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_8_fork (
    .io_input_valid          (signalInput_8_valid                               ), //i
    .io_input_ready          (signalInput_8_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_8_payload                             ), //i
    .io_outputs_0_valid      (signalInput_8_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_8_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_8_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_8_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_8_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_8_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_9_fork (
    .io_input_valid          (signalInput_9_valid                               ), //i
    .io_input_ready          (signalInput_9_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_9_payload                             ), //i
    .io_outputs_0_valid      (signalInput_9_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_9_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_9_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_9_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_9_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_9_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_10_fork (
    .io_input_valid          (signalInput_10_valid                               ), //i
    .io_input_ready          (signalInput_10_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_10_payload                             ), //i
    .io_outputs_0_valid      (signalInput_10_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_10_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_10_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_10_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_10_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_10_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_11_fork (
    .io_input_valid          (signalInput_11_valid                               ), //i
    .io_input_ready          (signalInput_11_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_11_payload                             ), //i
    .io_outputs_0_valid      (signalInput_11_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_11_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_11_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_11_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_11_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_11_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_12_fork (
    .io_input_valid          (signalInput_12_valid                               ), //i
    .io_input_ready          (signalInput_12_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_12_payload                             ), //i
    .io_outputs_0_valid      (signalInput_12_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_12_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_12_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_12_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_12_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_12_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_13_fork (
    .io_input_valid          (signalInput_13_valid                               ), //i
    .io_input_ready          (signalInput_13_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_13_payload                             ), //i
    .io_outputs_0_valid      (signalInput_13_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_13_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_13_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_13_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_13_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_13_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_14_fork (
    .io_input_valid          (signalInput_14_valid                               ), //i
    .io_input_ready          (signalInput_14_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_14_payload                             ), //i
    .io_outputs_0_valid      (signalInput_14_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_14_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_14_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_14_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_14_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_14_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_15_fork (
    .io_input_valid          (signalInput_15_valid                               ), //i
    .io_input_ready          (signalInput_15_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_15_payload                             ), //i
    .io_outputs_0_valid      (signalInput_15_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_15_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_15_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_15_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_15_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_15_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_16_fork (
    .io_input_valid          (signalInput_16_valid                               ), //i
    .io_input_ready          (signalInput_16_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_16_payload                             ), //i
    .io_outputs_0_valid      (signalInput_16_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_16_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_16_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_16_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_16_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_16_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_17_fork (
    .io_input_valid          (signalInput_17_valid                               ), //i
    .io_input_ready          (signalInput_17_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_17_payload                             ), //i
    .io_outputs_0_valid      (signalInput_17_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_17_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_17_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_17_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_17_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_17_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_18_fork (
    .io_input_valid          (signalInput_18_valid                               ), //i
    .io_input_ready          (signalInput_18_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_18_payload                             ), //i
    .io_outputs_0_valid      (signalInput_18_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_18_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_18_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_18_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_18_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_18_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_19_fork (
    .io_input_valid          (signalInput_19_valid                               ), //i
    .io_input_ready          (signalInput_19_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_19_payload                             ), //i
    .io_outputs_0_valid      (signalInput_19_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_19_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_19_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_19_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_19_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_19_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_20_fork (
    .io_input_valid          (signalInput_20_valid                               ), //i
    .io_input_ready          (signalInput_20_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_20_payload                             ), //i
    .io_outputs_0_valid      (signalInput_20_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_20_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_20_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_20_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_20_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_20_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_21_fork (
    .io_input_valid          (signalInput_21_valid                               ), //i
    .io_input_ready          (signalInput_21_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_21_payload                             ), //i
    .io_outputs_0_valid      (signalInput_21_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_21_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_21_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_21_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_21_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_21_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_22_fork (
    .io_input_valid          (signalInput_22_valid                               ), //i
    .io_input_ready          (signalInput_22_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_22_payload                             ), //i
    .io_outputs_0_valid      (signalInput_22_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_22_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_22_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_22_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_22_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_22_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_23_fork (
    .io_input_valid          (signalInput_23_valid                               ), //i
    .io_input_ready          (signalInput_23_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_23_payload                             ), //i
    .io_outputs_0_valid      (signalInput_23_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_23_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_23_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_23_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_23_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_23_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_24_fork (
    .io_input_valid          (signalInput_24_valid                               ), //i
    .io_input_ready          (signalInput_24_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_24_payload                             ), //i
    .io_outputs_0_valid      (signalInput_24_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_24_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_24_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_24_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_24_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_24_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_25_fork (
    .io_input_valid          (signalInput_25_valid                               ), //i
    .io_input_ready          (signalInput_25_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_25_payload                             ), //i
    .io_outputs_0_valid      (signalInput_25_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_25_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_25_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_25_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_25_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_25_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_26_fork (
    .io_input_valid          (signalInput_26_valid                               ), //i
    .io_input_ready          (signalInput_26_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_26_payload                             ), //i
    .io_outputs_0_valid      (signalInput_26_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_26_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_26_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_26_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_26_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_26_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_27_fork (
    .io_input_valid          (signalInput_27_valid                               ), //i
    .io_input_ready          (signalInput_27_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_27_payload                             ), //i
    .io_outputs_0_valid      (signalInput_27_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_27_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_27_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_27_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_27_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_27_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_28_fork (
    .io_input_valid          (signalInput_28_valid                               ), //i
    .io_input_ready          (signalInput_28_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_28_payload                             ), //i
    .io_outputs_0_valid      (signalInput_28_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_28_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_28_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_28_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_28_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_28_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_29_fork (
    .io_input_valid          (signalInput_29_valid                               ), //i
    .io_input_ready          (signalInput_29_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_29_payload                             ), //i
    .io_outputs_0_valid      (signalInput_29_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_29_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_29_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_29_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_29_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_29_fork_io_outputs_1_payload           )  //o
  );
  StreamFork signalInput_30_fork (
    .io_input_valid          (signalInput_30_valid                               ), //i
    .io_input_ready          (signalInput_30_fork_io_input_ready                 ), //o
    .io_input_payload        (signalInput_30_payload                             ), //i
    .io_outputs_0_valid      (signalInput_30_fork_io_outputs_0_valid             ), //o
    .io_outputs_0_ready      (signalInput_30_fork_io_outputs_0_ready             ), //i
    .io_outputs_0_payload    (signalInput_30_fork_io_outputs_0_payload           ), //o
    .io_outputs_1_valid      (signalInput_30_fork_io_outputs_1_valid             ), //o
    .io_outputs_1_ready      (signalInput_30_fork_io_outputs_1_translated_ready  ), //i
    .io_outputs_1_payload    (signalInput_30_fork_io_outputs_1_payload           )  //o
  );
  assign signalInput_0_ready = signalInput_0_fork_io_input_ready;
  always @(*) begin
    signalInput_0_fork_io_outputs_0_ready = signalInput_0_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342) begin
      signalInput_0_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! signalInput_0_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_0_fork_io_outputs_0_m2sPipe_valid = signalInput_0_fork_io_outputs_0_rValid;
  assign signalInput_0_fork_io_outputs_0_m2sPipe_payload = signalInput_0_fork_io_outputs_0_rData;
  assign signalInput_0_fork_io_outputs_1_translated_valid = signalInput_0_fork_io_outputs_1_valid;
  assign signalInput_0_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_0_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_0_fork_io_outputs_1_translated_payload};
  assign mulOut_0_valid = signalInput_0_fork_io_outputs_1_translated_valid;
  assign signalInput_0_fork_io_outputs_1_translated_ready = mulOut_0_ready;
  assign mulOut_0_payload = signalInput_0_fork_io_outputs_1_translated_payload;
  assign signalInput_1_ready = signalInput_1_fork_io_input_ready;
  always @(*) begin
    signalInput_1_fork_io_outputs_0_ready = signalInput_1_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      signalInput_1_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! signalInput_1_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_1_fork_io_outputs_0_m2sPipe_valid = signalInput_1_fork_io_outputs_0_rValid;
  assign signalInput_1_fork_io_outputs_0_m2sPipe_payload = signalInput_1_fork_io_outputs_0_rData;
  assign signalInput_1_fork_io_outputs_1_translated_valid = signalInput_1_fork_io_outputs_1_valid;
  assign signalInput_1_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_1_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_1_fork_io_outputs_1_translated_payload};
  assign mulOut_1_valid = signalInput_1_fork_io_outputs_1_translated_valid;
  assign signalInput_1_fork_io_outputs_1_translated_ready = mulOut_1_ready;
  assign mulOut_1_payload = signalInput_1_fork_io_outputs_1_translated_payload;
  assign signalInput_2_ready = signalInput_2_fork_io_input_ready;
  always @(*) begin
    signalInput_2_fork_io_outputs_0_ready = signalInput_2_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      signalInput_2_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! signalInput_2_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_2_fork_io_outputs_0_m2sPipe_valid = signalInput_2_fork_io_outputs_0_rValid;
  assign signalInput_2_fork_io_outputs_0_m2sPipe_payload = signalInput_2_fork_io_outputs_0_rData;
  assign signalInput_2_fork_io_outputs_1_translated_valid = signalInput_2_fork_io_outputs_1_valid;
  assign signalInput_2_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_2_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_2_fork_io_outputs_1_translated_payload};
  assign mulOut_2_valid = signalInput_2_fork_io_outputs_1_translated_valid;
  assign signalInput_2_fork_io_outputs_1_translated_ready = mulOut_2_ready;
  assign mulOut_2_payload = signalInput_2_fork_io_outputs_1_translated_payload;
  assign signalInput_3_ready = signalInput_3_fork_io_input_ready;
  always @(*) begin
    signalInput_3_fork_io_outputs_0_ready = signalInput_3_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_3) begin
      signalInput_3_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! signalInput_3_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_3_fork_io_outputs_0_m2sPipe_valid = signalInput_3_fork_io_outputs_0_rValid;
  assign signalInput_3_fork_io_outputs_0_m2sPipe_payload = signalInput_3_fork_io_outputs_0_rData;
  assign signalInput_3_fork_io_outputs_1_translated_valid = signalInput_3_fork_io_outputs_1_valid;
  assign signalInput_3_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_3_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_3_fork_io_outputs_1_translated_payload};
  assign mulOut_3_valid = signalInput_3_fork_io_outputs_1_translated_valid;
  assign signalInput_3_fork_io_outputs_1_translated_ready = mulOut_3_ready;
  assign mulOut_3_payload = signalInput_3_fork_io_outputs_1_translated_payload;
  assign signalInput_4_ready = signalInput_4_fork_io_input_ready;
  always @(*) begin
    signalInput_4_fork_io_outputs_0_ready = signalInput_4_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_4) begin
      signalInput_4_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! signalInput_4_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_4_fork_io_outputs_0_m2sPipe_valid = signalInput_4_fork_io_outputs_0_rValid;
  assign signalInput_4_fork_io_outputs_0_m2sPipe_payload = signalInput_4_fork_io_outputs_0_rData;
  assign signalInput_4_fork_io_outputs_1_translated_valid = signalInput_4_fork_io_outputs_1_valid;
  assign signalInput_4_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_4_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_4_fork_io_outputs_1_translated_payload};
  assign mulOut_4_valid = signalInput_4_fork_io_outputs_1_translated_valid;
  assign signalInput_4_fork_io_outputs_1_translated_ready = mulOut_4_ready;
  assign mulOut_4_payload = signalInput_4_fork_io_outputs_1_translated_payload;
  assign signalInput_5_ready = signalInput_5_fork_io_input_ready;
  always @(*) begin
    signalInput_5_fork_io_outputs_0_ready = signalInput_5_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_5) begin
      signalInput_5_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! signalInput_5_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_5_fork_io_outputs_0_m2sPipe_valid = signalInput_5_fork_io_outputs_0_rValid;
  assign signalInput_5_fork_io_outputs_0_m2sPipe_payload = signalInput_5_fork_io_outputs_0_rData;
  assign signalInput_5_fork_io_outputs_1_translated_valid = signalInput_5_fork_io_outputs_1_valid;
  assign signalInput_5_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_5_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_5_fork_io_outputs_1_translated_payload};
  assign mulOut_5_valid = signalInput_5_fork_io_outputs_1_translated_valid;
  assign signalInput_5_fork_io_outputs_1_translated_ready = mulOut_5_ready;
  assign mulOut_5_payload = signalInput_5_fork_io_outputs_1_translated_payload;
  assign signalInput_6_ready = signalInput_6_fork_io_input_ready;
  always @(*) begin
    signalInput_6_fork_io_outputs_0_ready = signalInput_6_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_6) begin
      signalInput_6_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_6 = (! signalInput_6_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_6_fork_io_outputs_0_m2sPipe_valid = signalInput_6_fork_io_outputs_0_rValid;
  assign signalInput_6_fork_io_outputs_0_m2sPipe_payload = signalInput_6_fork_io_outputs_0_rData;
  assign signalInput_6_fork_io_outputs_1_translated_valid = signalInput_6_fork_io_outputs_1_valid;
  assign signalInput_6_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_6_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_6_fork_io_outputs_1_translated_payload};
  assign mulOut_6_valid = signalInput_6_fork_io_outputs_1_translated_valid;
  assign signalInput_6_fork_io_outputs_1_translated_ready = mulOut_6_ready;
  assign mulOut_6_payload = signalInput_6_fork_io_outputs_1_translated_payload;
  assign signalInput_7_ready = signalInput_7_fork_io_input_ready;
  always @(*) begin
    signalInput_7_fork_io_outputs_0_ready = signalInput_7_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_7) begin
      signalInput_7_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_7 = (! signalInput_7_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_7_fork_io_outputs_0_m2sPipe_valid = signalInput_7_fork_io_outputs_0_rValid;
  assign signalInput_7_fork_io_outputs_0_m2sPipe_payload = signalInput_7_fork_io_outputs_0_rData;
  assign signalInput_7_fork_io_outputs_1_translated_valid = signalInput_7_fork_io_outputs_1_valid;
  assign signalInput_7_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_7_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_7_fork_io_outputs_1_translated_payload};
  assign mulOut_7_valid = signalInput_7_fork_io_outputs_1_translated_valid;
  assign signalInput_7_fork_io_outputs_1_translated_ready = mulOut_7_ready;
  assign mulOut_7_payload = signalInput_7_fork_io_outputs_1_translated_payload;
  assign signalInput_8_ready = signalInput_8_fork_io_input_ready;
  always @(*) begin
    signalInput_8_fork_io_outputs_0_ready = signalInput_8_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_8) begin
      signalInput_8_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_8 = (! signalInput_8_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_8_fork_io_outputs_0_m2sPipe_valid = signalInput_8_fork_io_outputs_0_rValid;
  assign signalInput_8_fork_io_outputs_0_m2sPipe_payload = signalInput_8_fork_io_outputs_0_rData;
  assign signalInput_8_fork_io_outputs_1_translated_valid = signalInput_8_fork_io_outputs_1_valid;
  assign signalInput_8_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_8_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_8_fork_io_outputs_1_translated_payload};
  assign mulOut_8_valid = signalInput_8_fork_io_outputs_1_translated_valid;
  assign signalInput_8_fork_io_outputs_1_translated_ready = mulOut_8_ready;
  assign mulOut_8_payload = signalInput_8_fork_io_outputs_1_translated_payload;
  assign signalInput_9_ready = signalInput_9_fork_io_input_ready;
  always @(*) begin
    signalInput_9_fork_io_outputs_0_ready = signalInput_9_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_9) begin
      signalInput_9_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_9 = (! signalInput_9_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_9_fork_io_outputs_0_m2sPipe_valid = signalInput_9_fork_io_outputs_0_rValid;
  assign signalInput_9_fork_io_outputs_0_m2sPipe_payload = signalInput_9_fork_io_outputs_0_rData;
  assign signalInput_9_fork_io_outputs_1_translated_valid = signalInput_9_fork_io_outputs_1_valid;
  assign signalInput_9_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_9_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_9_fork_io_outputs_1_translated_payload};
  assign mulOut_9_valid = signalInput_9_fork_io_outputs_1_translated_valid;
  assign signalInput_9_fork_io_outputs_1_translated_ready = mulOut_9_ready;
  assign mulOut_9_payload = signalInput_9_fork_io_outputs_1_translated_payload;
  assign signalInput_10_ready = signalInput_10_fork_io_input_ready;
  always @(*) begin
    signalInput_10_fork_io_outputs_0_ready = signalInput_10_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_10) begin
      signalInput_10_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_10 = (! signalInput_10_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_10_fork_io_outputs_0_m2sPipe_valid = signalInput_10_fork_io_outputs_0_rValid;
  assign signalInput_10_fork_io_outputs_0_m2sPipe_payload = signalInput_10_fork_io_outputs_0_rData;
  assign signalInput_10_fork_io_outputs_1_translated_valid = signalInput_10_fork_io_outputs_1_valid;
  assign signalInput_10_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_10_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_10_fork_io_outputs_1_translated_payload};
  assign mulOut_10_valid = signalInput_10_fork_io_outputs_1_translated_valid;
  assign signalInput_10_fork_io_outputs_1_translated_ready = mulOut_10_ready;
  assign mulOut_10_payload = signalInput_10_fork_io_outputs_1_translated_payload;
  assign signalInput_11_ready = signalInput_11_fork_io_input_ready;
  always @(*) begin
    signalInput_11_fork_io_outputs_0_ready = signalInput_11_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_11) begin
      signalInput_11_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_11 = (! signalInput_11_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_11_fork_io_outputs_0_m2sPipe_valid = signalInput_11_fork_io_outputs_0_rValid;
  assign signalInput_11_fork_io_outputs_0_m2sPipe_payload = signalInput_11_fork_io_outputs_0_rData;
  assign signalInput_11_fork_io_outputs_1_translated_valid = signalInput_11_fork_io_outputs_1_valid;
  assign signalInput_11_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_11_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_11_fork_io_outputs_1_translated_payload};
  assign mulOut_11_valid = signalInput_11_fork_io_outputs_1_translated_valid;
  assign signalInput_11_fork_io_outputs_1_translated_ready = mulOut_11_ready;
  assign mulOut_11_payload = signalInput_11_fork_io_outputs_1_translated_payload;
  assign signalInput_12_ready = signalInput_12_fork_io_input_ready;
  always @(*) begin
    signalInput_12_fork_io_outputs_0_ready = signalInput_12_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_12) begin
      signalInput_12_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_12 = (! signalInput_12_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_12_fork_io_outputs_0_m2sPipe_valid = signalInput_12_fork_io_outputs_0_rValid;
  assign signalInput_12_fork_io_outputs_0_m2sPipe_payload = signalInput_12_fork_io_outputs_0_rData;
  assign signalInput_12_fork_io_outputs_1_translated_valid = signalInput_12_fork_io_outputs_1_valid;
  assign signalInput_12_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_12_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_12_fork_io_outputs_1_translated_payload};
  assign mulOut_12_valid = signalInput_12_fork_io_outputs_1_translated_valid;
  assign signalInput_12_fork_io_outputs_1_translated_ready = mulOut_12_ready;
  assign mulOut_12_payload = signalInput_12_fork_io_outputs_1_translated_payload;
  assign signalInput_13_ready = signalInput_13_fork_io_input_ready;
  always @(*) begin
    signalInput_13_fork_io_outputs_0_ready = signalInput_13_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_13) begin
      signalInput_13_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_13 = (! signalInput_13_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_13_fork_io_outputs_0_m2sPipe_valid = signalInput_13_fork_io_outputs_0_rValid;
  assign signalInput_13_fork_io_outputs_0_m2sPipe_payload = signalInput_13_fork_io_outputs_0_rData;
  assign signalInput_13_fork_io_outputs_1_translated_valid = signalInput_13_fork_io_outputs_1_valid;
  assign signalInput_13_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_13_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_13_fork_io_outputs_1_translated_payload};
  assign mulOut_13_valid = signalInput_13_fork_io_outputs_1_translated_valid;
  assign signalInput_13_fork_io_outputs_1_translated_ready = mulOut_13_ready;
  assign mulOut_13_payload = signalInput_13_fork_io_outputs_1_translated_payload;
  assign signalInput_14_ready = signalInput_14_fork_io_input_ready;
  always @(*) begin
    signalInput_14_fork_io_outputs_0_ready = signalInput_14_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_14) begin
      signalInput_14_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_14 = (! signalInput_14_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_14_fork_io_outputs_0_m2sPipe_valid = signalInput_14_fork_io_outputs_0_rValid;
  assign signalInput_14_fork_io_outputs_0_m2sPipe_payload = signalInput_14_fork_io_outputs_0_rData;
  assign signalInput_14_fork_io_outputs_1_translated_valid = signalInput_14_fork_io_outputs_1_valid;
  assign signalInput_14_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_14_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_14_fork_io_outputs_1_translated_payload};
  assign mulOut_14_valid = signalInput_14_fork_io_outputs_1_translated_valid;
  assign signalInput_14_fork_io_outputs_1_translated_ready = mulOut_14_ready;
  assign mulOut_14_payload = signalInput_14_fork_io_outputs_1_translated_payload;
  assign signalInput_15_ready = signalInput_15_fork_io_input_ready;
  always @(*) begin
    signalInput_15_fork_io_outputs_0_ready = signalInput_15_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_15) begin
      signalInput_15_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_15 = (! signalInput_15_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_15_fork_io_outputs_0_m2sPipe_valid = signalInput_15_fork_io_outputs_0_rValid;
  assign signalInput_15_fork_io_outputs_0_m2sPipe_payload = signalInput_15_fork_io_outputs_0_rData;
  assign signalInput_15_fork_io_outputs_1_translated_valid = signalInput_15_fork_io_outputs_1_valid;
  assign signalInput_15_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_15_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_15_fork_io_outputs_1_translated_payload};
  assign mulOut_15_valid = signalInput_15_fork_io_outputs_1_translated_valid;
  assign signalInput_15_fork_io_outputs_1_translated_ready = mulOut_15_ready;
  assign mulOut_15_payload = signalInput_15_fork_io_outputs_1_translated_payload;
  assign signalInput_16_ready = signalInput_16_fork_io_input_ready;
  always @(*) begin
    signalInput_16_fork_io_outputs_0_ready = signalInput_16_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_16) begin
      signalInput_16_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_16 = (! signalInput_16_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_16_fork_io_outputs_0_m2sPipe_valid = signalInput_16_fork_io_outputs_0_rValid;
  assign signalInput_16_fork_io_outputs_0_m2sPipe_payload = signalInput_16_fork_io_outputs_0_rData;
  assign signalInput_16_fork_io_outputs_1_translated_valid = signalInput_16_fork_io_outputs_1_valid;
  assign signalInput_16_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_16_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_16_fork_io_outputs_1_translated_payload};
  assign mulOut_16_valid = signalInput_16_fork_io_outputs_1_translated_valid;
  assign signalInput_16_fork_io_outputs_1_translated_ready = mulOut_16_ready;
  assign mulOut_16_payload = signalInput_16_fork_io_outputs_1_translated_payload;
  assign signalInput_17_ready = signalInput_17_fork_io_input_ready;
  always @(*) begin
    signalInput_17_fork_io_outputs_0_ready = signalInput_17_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_17) begin
      signalInput_17_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_17 = (! signalInput_17_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_17_fork_io_outputs_0_m2sPipe_valid = signalInput_17_fork_io_outputs_0_rValid;
  assign signalInput_17_fork_io_outputs_0_m2sPipe_payload = signalInput_17_fork_io_outputs_0_rData;
  assign signalInput_17_fork_io_outputs_1_translated_valid = signalInput_17_fork_io_outputs_1_valid;
  assign signalInput_17_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_17_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_17_fork_io_outputs_1_translated_payload};
  assign mulOut_17_valid = signalInput_17_fork_io_outputs_1_translated_valid;
  assign signalInput_17_fork_io_outputs_1_translated_ready = mulOut_17_ready;
  assign mulOut_17_payload = signalInput_17_fork_io_outputs_1_translated_payload;
  assign signalInput_18_ready = signalInput_18_fork_io_input_ready;
  always @(*) begin
    signalInput_18_fork_io_outputs_0_ready = signalInput_18_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_18) begin
      signalInput_18_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_18 = (! signalInput_18_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_18_fork_io_outputs_0_m2sPipe_valid = signalInput_18_fork_io_outputs_0_rValid;
  assign signalInput_18_fork_io_outputs_0_m2sPipe_payload = signalInput_18_fork_io_outputs_0_rData;
  assign signalInput_18_fork_io_outputs_1_translated_valid = signalInput_18_fork_io_outputs_1_valid;
  assign signalInput_18_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_18_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_18_fork_io_outputs_1_translated_payload};
  assign mulOut_18_valid = signalInput_18_fork_io_outputs_1_translated_valid;
  assign signalInput_18_fork_io_outputs_1_translated_ready = mulOut_18_ready;
  assign mulOut_18_payload = signalInput_18_fork_io_outputs_1_translated_payload;
  assign signalInput_19_ready = signalInput_19_fork_io_input_ready;
  always @(*) begin
    signalInput_19_fork_io_outputs_0_ready = signalInput_19_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_19) begin
      signalInput_19_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_19 = (! signalInput_19_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_19_fork_io_outputs_0_m2sPipe_valid = signalInput_19_fork_io_outputs_0_rValid;
  assign signalInput_19_fork_io_outputs_0_m2sPipe_payload = signalInput_19_fork_io_outputs_0_rData;
  assign signalInput_19_fork_io_outputs_1_translated_valid = signalInput_19_fork_io_outputs_1_valid;
  assign signalInput_19_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_19_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_19_fork_io_outputs_1_translated_payload};
  assign mulOut_19_valid = signalInput_19_fork_io_outputs_1_translated_valid;
  assign signalInput_19_fork_io_outputs_1_translated_ready = mulOut_19_ready;
  assign mulOut_19_payload = signalInput_19_fork_io_outputs_1_translated_payload;
  assign signalInput_20_ready = signalInput_20_fork_io_input_ready;
  always @(*) begin
    signalInput_20_fork_io_outputs_0_ready = signalInput_20_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_20) begin
      signalInput_20_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_20 = (! signalInput_20_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_20_fork_io_outputs_0_m2sPipe_valid = signalInput_20_fork_io_outputs_0_rValid;
  assign signalInput_20_fork_io_outputs_0_m2sPipe_payload = signalInput_20_fork_io_outputs_0_rData;
  assign signalInput_20_fork_io_outputs_1_translated_valid = signalInput_20_fork_io_outputs_1_valid;
  assign signalInput_20_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_20_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_20_fork_io_outputs_1_translated_payload};
  assign mulOut_20_valid = signalInput_20_fork_io_outputs_1_translated_valid;
  assign signalInput_20_fork_io_outputs_1_translated_ready = mulOut_20_ready;
  assign mulOut_20_payload = signalInput_20_fork_io_outputs_1_translated_payload;
  assign signalInput_21_ready = signalInput_21_fork_io_input_ready;
  always @(*) begin
    signalInput_21_fork_io_outputs_0_ready = signalInput_21_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_21) begin
      signalInput_21_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_21 = (! signalInput_21_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_21_fork_io_outputs_0_m2sPipe_valid = signalInput_21_fork_io_outputs_0_rValid;
  assign signalInput_21_fork_io_outputs_0_m2sPipe_payload = signalInput_21_fork_io_outputs_0_rData;
  assign signalInput_21_fork_io_outputs_1_translated_valid = signalInput_21_fork_io_outputs_1_valid;
  assign signalInput_21_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_21_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_21_fork_io_outputs_1_translated_payload};
  assign mulOut_21_valid = signalInput_21_fork_io_outputs_1_translated_valid;
  assign signalInput_21_fork_io_outputs_1_translated_ready = mulOut_21_ready;
  assign mulOut_21_payload = signalInput_21_fork_io_outputs_1_translated_payload;
  assign signalInput_22_ready = signalInput_22_fork_io_input_ready;
  always @(*) begin
    signalInput_22_fork_io_outputs_0_ready = signalInput_22_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_22) begin
      signalInput_22_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_22 = (! signalInput_22_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_22_fork_io_outputs_0_m2sPipe_valid = signalInput_22_fork_io_outputs_0_rValid;
  assign signalInput_22_fork_io_outputs_0_m2sPipe_payload = signalInput_22_fork_io_outputs_0_rData;
  assign signalInput_22_fork_io_outputs_1_translated_valid = signalInput_22_fork_io_outputs_1_valid;
  assign signalInput_22_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_22_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_22_fork_io_outputs_1_translated_payload};
  assign mulOut_22_valid = signalInput_22_fork_io_outputs_1_translated_valid;
  assign signalInput_22_fork_io_outputs_1_translated_ready = mulOut_22_ready;
  assign mulOut_22_payload = signalInput_22_fork_io_outputs_1_translated_payload;
  assign signalInput_23_ready = signalInput_23_fork_io_input_ready;
  always @(*) begin
    signalInput_23_fork_io_outputs_0_ready = signalInput_23_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_23) begin
      signalInput_23_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_23 = (! signalInput_23_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_23_fork_io_outputs_0_m2sPipe_valid = signalInput_23_fork_io_outputs_0_rValid;
  assign signalInput_23_fork_io_outputs_0_m2sPipe_payload = signalInput_23_fork_io_outputs_0_rData;
  assign signalInput_23_fork_io_outputs_1_translated_valid = signalInput_23_fork_io_outputs_1_valid;
  assign signalInput_23_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_23_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_23_fork_io_outputs_1_translated_payload};
  assign mulOut_23_valid = signalInput_23_fork_io_outputs_1_translated_valid;
  assign signalInput_23_fork_io_outputs_1_translated_ready = mulOut_23_ready;
  assign mulOut_23_payload = signalInput_23_fork_io_outputs_1_translated_payload;
  assign signalInput_24_ready = signalInput_24_fork_io_input_ready;
  always @(*) begin
    signalInput_24_fork_io_outputs_0_ready = signalInput_24_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_24) begin
      signalInput_24_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_24 = (! signalInput_24_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_24_fork_io_outputs_0_m2sPipe_valid = signalInput_24_fork_io_outputs_0_rValid;
  assign signalInput_24_fork_io_outputs_0_m2sPipe_payload = signalInput_24_fork_io_outputs_0_rData;
  assign signalInput_24_fork_io_outputs_1_translated_valid = signalInput_24_fork_io_outputs_1_valid;
  assign signalInput_24_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_24_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_24_fork_io_outputs_1_translated_payload};
  assign mulOut_24_valid = signalInput_24_fork_io_outputs_1_translated_valid;
  assign signalInput_24_fork_io_outputs_1_translated_ready = mulOut_24_ready;
  assign mulOut_24_payload = signalInput_24_fork_io_outputs_1_translated_payload;
  assign signalInput_25_ready = signalInput_25_fork_io_input_ready;
  always @(*) begin
    signalInput_25_fork_io_outputs_0_ready = signalInput_25_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_25) begin
      signalInput_25_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_25 = (! signalInput_25_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_25_fork_io_outputs_0_m2sPipe_valid = signalInput_25_fork_io_outputs_0_rValid;
  assign signalInput_25_fork_io_outputs_0_m2sPipe_payload = signalInput_25_fork_io_outputs_0_rData;
  assign signalInput_25_fork_io_outputs_1_translated_valid = signalInput_25_fork_io_outputs_1_valid;
  assign signalInput_25_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_25_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_25_fork_io_outputs_1_translated_payload};
  assign mulOut_25_valid = signalInput_25_fork_io_outputs_1_translated_valid;
  assign signalInput_25_fork_io_outputs_1_translated_ready = mulOut_25_ready;
  assign mulOut_25_payload = signalInput_25_fork_io_outputs_1_translated_payload;
  assign signalInput_26_ready = signalInput_26_fork_io_input_ready;
  always @(*) begin
    signalInput_26_fork_io_outputs_0_ready = signalInput_26_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_26) begin
      signalInput_26_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_26 = (! signalInput_26_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_26_fork_io_outputs_0_m2sPipe_valid = signalInput_26_fork_io_outputs_0_rValid;
  assign signalInput_26_fork_io_outputs_0_m2sPipe_payload = signalInput_26_fork_io_outputs_0_rData;
  assign signalInput_26_fork_io_outputs_1_translated_valid = signalInput_26_fork_io_outputs_1_valid;
  assign signalInput_26_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_26_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_26_fork_io_outputs_1_translated_payload};
  assign mulOut_26_valid = signalInput_26_fork_io_outputs_1_translated_valid;
  assign signalInput_26_fork_io_outputs_1_translated_ready = mulOut_26_ready;
  assign mulOut_26_payload = signalInput_26_fork_io_outputs_1_translated_payload;
  assign signalInput_27_ready = signalInput_27_fork_io_input_ready;
  always @(*) begin
    signalInput_27_fork_io_outputs_0_ready = signalInput_27_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_27) begin
      signalInput_27_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_27 = (! signalInput_27_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_27_fork_io_outputs_0_m2sPipe_valid = signalInput_27_fork_io_outputs_0_rValid;
  assign signalInput_27_fork_io_outputs_0_m2sPipe_payload = signalInput_27_fork_io_outputs_0_rData;
  assign signalInput_27_fork_io_outputs_1_translated_valid = signalInput_27_fork_io_outputs_1_valid;
  assign signalInput_27_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_27_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_27_fork_io_outputs_1_translated_payload};
  assign mulOut_27_valid = signalInput_27_fork_io_outputs_1_translated_valid;
  assign signalInput_27_fork_io_outputs_1_translated_ready = mulOut_27_ready;
  assign mulOut_27_payload = signalInput_27_fork_io_outputs_1_translated_payload;
  assign signalInput_28_ready = signalInput_28_fork_io_input_ready;
  always @(*) begin
    signalInput_28_fork_io_outputs_0_ready = signalInput_28_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_28) begin
      signalInput_28_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_28 = (! signalInput_28_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_28_fork_io_outputs_0_m2sPipe_valid = signalInput_28_fork_io_outputs_0_rValid;
  assign signalInput_28_fork_io_outputs_0_m2sPipe_payload = signalInput_28_fork_io_outputs_0_rData;
  assign signalInput_28_fork_io_outputs_1_translated_valid = signalInput_28_fork_io_outputs_1_valid;
  assign signalInput_28_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_28_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_28_fork_io_outputs_1_translated_payload};
  assign mulOut_28_valid = signalInput_28_fork_io_outputs_1_translated_valid;
  assign signalInput_28_fork_io_outputs_1_translated_ready = mulOut_28_ready;
  assign mulOut_28_payload = signalInput_28_fork_io_outputs_1_translated_payload;
  assign signalInput_29_ready = signalInput_29_fork_io_input_ready;
  always @(*) begin
    signalInput_29_fork_io_outputs_0_ready = signalInput_29_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_29) begin
      signalInput_29_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_29 = (! signalInput_29_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_29_fork_io_outputs_0_m2sPipe_valid = signalInput_29_fork_io_outputs_0_rValid;
  assign signalInput_29_fork_io_outputs_0_m2sPipe_payload = signalInput_29_fork_io_outputs_0_rData;
  assign signalInput_29_fork_io_outputs_1_translated_valid = signalInput_29_fork_io_outputs_1_valid;
  assign signalInput_29_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_29_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_29_fork_io_outputs_1_translated_payload};
  assign mulOut_29_valid = signalInput_29_fork_io_outputs_1_translated_valid;
  assign signalInput_29_fork_io_outputs_1_translated_ready = mulOut_29_ready;
  assign mulOut_29_payload = signalInput_29_fork_io_outputs_1_translated_payload;
  assign signalInput_30_ready = signalInput_30_fork_io_input_ready;
  always @(*) begin
    signalInput_30_fork_io_outputs_0_ready = signalInput_30_fork_io_outputs_0_m2sPipe_ready;
    if(when_Stream_l342_30) begin
      signalInput_30_fork_io_outputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_30 = (! signalInput_30_fork_io_outputs_0_m2sPipe_valid);
  assign signalInput_30_fork_io_outputs_0_m2sPipe_valid = signalInput_30_fork_io_outputs_0_rValid;
  assign signalInput_30_fork_io_outputs_0_m2sPipe_payload = signalInput_30_fork_io_outputs_0_rData;
  assign signalInput_30_fork_io_outputs_1_translated_valid = signalInput_30_fork_io_outputs_1_valid;
  assign signalInput_30_fork_io_outputs_1_translated_payload = {{3{_zz_signalInput_30_fork_io_outputs_1_translated_payload[16]}}, _zz_signalInput_30_fork_io_outputs_1_translated_payload};
  assign mulOut_30_valid = signalInput_30_fork_io_outputs_1_translated_valid;
  assign signalInput_30_fork_io_outputs_1_translated_ready = mulOut_30_ready;
  assign mulOut_30_payload = signalInput_30_fork_io_outputs_1_translated_payload;
  assign signalInput_0_valid = io_input_valid;
  assign io_input_ready = signalInput_0_ready;
  assign signalInput_0_payload = io_input_payload;
  assign signalInput_1_valid = signalInput_0_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_0_fork_io_outputs_0_m2sPipe_ready = signalInput_1_ready;
  assign signalInput_1_payload = signalInput_0_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_2_valid = signalInput_1_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_1_fork_io_outputs_0_m2sPipe_ready = signalInput_2_ready;
  assign signalInput_2_payload = signalInput_1_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_3_valid = signalInput_2_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_2_fork_io_outputs_0_m2sPipe_ready = signalInput_3_ready;
  assign signalInput_3_payload = signalInput_2_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_4_valid = signalInput_3_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_3_fork_io_outputs_0_m2sPipe_ready = signalInput_4_ready;
  assign signalInput_4_payload = signalInput_3_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_5_valid = signalInput_4_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_4_fork_io_outputs_0_m2sPipe_ready = signalInput_5_ready;
  assign signalInput_5_payload = signalInput_4_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_6_valid = signalInput_5_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_5_fork_io_outputs_0_m2sPipe_ready = signalInput_6_ready;
  assign signalInput_6_payload = signalInput_5_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_7_valid = signalInput_6_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_6_fork_io_outputs_0_m2sPipe_ready = signalInput_7_ready;
  assign signalInput_7_payload = signalInput_6_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_8_valid = signalInput_7_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_7_fork_io_outputs_0_m2sPipe_ready = signalInput_8_ready;
  assign signalInput_8_payload = signalInput_7_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_9_valid = signalInput_8_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_8_fork_io_outputs_0_m2sPipe_ready = signalInput_9_ready;
  assign signalInput_9_payload = signalInput_8_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_10_valid = signalInput_9_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_9_fork_io_outputs_0_m2sPipe_ready = signalInput_10_ready;
  assign signalInput_10_payload = signalInput_9_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_11_valid = signalInput_10_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_10_fork_io_outputs_0_m2sPipe_ready = signalInput_11_ready;
  assign signalInput_11_payload = signalInput_10_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_12_valid = signalInput_11_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_11_fork_io_outputs_0_m2sPipe_ready = signalInput_12_ready;
  assign signalInput_12_payload = signalInput_11_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_13_valid = signalInput_12_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_12_fork_io_outputs_0_m2sPipe_ready = signalInput_13_ready;
  assign signalInput_13_payload = signalInput_12_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_14_valid = signalInput_13_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_13_fork_io_outputs_0_m2sPipe_ready = signalInput_14_ready;
  assign signalInput_14_payload = signalInput_13_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_15_valid = signalInput_14_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_14_fork_io_outputs_0_m2sPipe_ready = signalInput_15_ready;
  assign signalInput_15_payload = signalInput_14_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_16_valid = signalInput_15_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_15_fork_io_outputs_0_m2sPipe_ready = signalInput_16_ready;
  assign signalInput_16_payload = signalInput_15_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_17_valid = signalInput_16_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_16_fork_io_outputs_0_m2sPipe_ready = signalInput_17_ready;
  assign signalInput_17_payload = signalInput_16_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_18_valid = signalInput_17_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_17_fork_io_outputs_0_m2sPipe_ready = signalInput_18_ready;
  assign signalInput_18_payload = signalInput_17_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_19_valid = signalInput_18_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_18_fork_io_outputs_0_m2sPipe_ready = signalInput_19_ready;
  assign signalInput_19_payload = signalInput_18_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_20_valid = signalInput_19_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_19_fork_io_outputs_0_m2sPipe_ready = signalInput_20_ready;
  assign signalInput_20_payload = signalInput_19_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_21_valid = signalInput_20_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_20_fork_io_outputs_0_m2sPipe_ready = signalInput_21_ready;
  assign signalInput_21_payload = signalInput_20_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_22_valid = signalInput_21_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_21_fork_io_outputs_0_m2sPipe_ready = signalInput_22_ready;
  assign signalInput_22_payload = signalInput_21_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_23_valid = signalInput_22_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_22_fork_io_outputs_0_m2sPipe_ready = signalInput_23_ready;
  assign signalInput_23_payload = signalInput_22_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_24_valid = signalInput_23_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_23_fork_io_outputs_0_m2sPipe_ready = signalInput_24_ready;
  assign signalInput_24_payload = signalInput_23_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_25_valid = signalInput_24_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_24_fork_io_outputs_0_m2sPipe_ready = signalInput_25_ready;
  assign signalInput_25_payload = signalInput_24_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_26_valid = signalInput_25_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_25_fork_io_outputs_0_m2sPipe_ready = signalInput_26_ready;
  assign signalInput_26_payload = signalInput_25_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_27_valid = signalInput_26_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_26_fork_io_outputs_0_m2sPipe_ready = signalInput_27_ready;
  assign signalInput_27_payload = signalInput_26_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_28_valid = signalInput_27_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_27_fork_io_outputs_0_m2sPipe_ready = signalInput_28_ready;
  assign signalInput_28_payload = signalInput_27_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_29_valid = signalInput_28_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_28_fork_io_outputs_0_m2sPipe_ready = signalInput_29_ready;
  assign signalInput_29_payload = signalInput_28_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_30_valid = signalInput_29_fork_io_outputs_0_m2sPipe_valid;
  assign signalInput_29_fork_io_outputs_0_m2sPipe_ready = signalInput_30_ready;
  assign signalInput_30_payload = signalInput_29_fork_io_outputs_0_m2sPipe_payload;
  assign signalInput_30_fork_io_outputs_0_m2sPipe_ready = 1'b1;
  assign io_multiplyResult_valid = ((((((((((((((((_zz_io_multiplyResult_valid && mulOut_15_valid) && mulOut_16_valid) && mulOut_17_valid) && mulOut_18_valid) && mulOut_19_valid) && mulOut_20_valid) && mulOut_21_valid) && mulOut_22_valid) && mulOut_23_valid) && mulOut_24_valid) && mulOut_25_valid) && mulOut_26_valid) && mulOut_27_valid) && mulOut_28_valid) && mulOut_29_valid) && mulOut_30_valid);
  assign mulOut_0_ready = io_multiplyResult_ready;
  assign mulOut_1_ready = io_multiplyResult_ready;
  assign mulOut_2_ready = io_multiplyResult_ready;
  assign mulOut_3_ready = io_multiplyResult_ready;
  assign mulOut_4_ready = io_multiplyResult_ready;
  assign mulOut_5_ready = io_multiplyResult_ready;
  assign mulOut_6_ready = io_multiplyResult_ready;
  assign mulOut_7_ready = io_multiplyResult_ready;
  assign mulOut_8_ready = io_multiplyResult_ready;
  assign mulOut_9_ready = io_multiplyResult_ready;
  assign mulOut_10_ready = io_multiplyResult_ready;
  assign mulOut_11_ready = io_multiplyResult_ready;
  assign mulOut_12_ready = io_multiplyResult_ready;
  assign mulOut_13_ready = io_multiplyResult_ready;
  assign mulOut_14_ready = io_multiplyResult_ready;
  assign mulOut_15_ready = io_multiplyResult_ready;
  assign mulOut_16_ready = io_multiplyResult_ready;
  assign mulOut_17_ready = io_multiplyResult_ready;
  assign mulOut_18_ready = io_multiplyResult_ready;
  assign mulOut_19_ready = io_multiplyResult_ready;
  assign mulOut_20_ready = io_multiplyResult_ready;
  assign mulOut_21_ready = io_multiplyResult_ready;
  assign mulOut_22_ready = io_multiplyResult_ready;
  assign mulOut_23_ready = io_multiplyResult_ready;
  assign mulOut_24_ready = io_multiplyResult_ready;
  assign mulOut_25_ready = io_multiplyResult_ready;
  assign mulOut_26_ready = io_multiplyResult_ready;
  assign mulOut_27_ready = io_multiplyResult_ready;
  assign mulOut_28_ready = io_multiplyResult_ready;
  assign mulOut_29_ready = io_multiplyResult_ready;
  assign mulOut_30_ready = io_multiplyResult_ready;
  assign io_multiplyResult_payload_0 = mulOut_0_payload;
  assign io_multiplyResult_payload_1 = mulOut_1_payload;
  assign io_multiplyResult_payload_2 = mulOut_2_payload;
  assign io_multiplyResult_payload_3 = mulOut_3_payload;
  assign io_multiplyResult_payload_4 = mulOut_4_payload;
  assign io_multiplyResult_payload_5 = mulOut_5_payload;
  assign io_multiplyResult_payload_6 = mulOut_6_payload;
  assign io_multiplyResult_payload_7 = mulOut_7_payload;
  assign io_multiplyResult_payload_8 = mulOut_8_payload;
  assign io_multiplyResult_payload_9 = mulOut_9_payload;
  assign io_multiplyResult_payload_10 = mulOut_10_payload;
  assign io_multiplyResult_payload_11 = mulOut_11_payload;
  assign io_multiplyResult_payload_12 = mulOut_12_payload;
  assign io_multiplyResult_payload_13 = mulOut_13_payload;
  assign io_multiplyResult_payload_14 = mulOut_14_payload;
  assign io_multiplyResult_payload_15 = mulOut_15_payload;
  assign io_multiplyResult_payload_16 = mulOut_16_payload;
  assign io_multiplyResult_payload_17 = mulOut_17_payload;
  assign io_multiplyResult_payload_18 = mulOut_18_payload;
  assign io_multiplyResult_payload_19 = mulOut_19_payload;
  assign io_multiplyResult_payload_20 = mulOut_20_payload;
  assign io_multiplyResult_payload_21 = mulOut_21_payload;
  assign io_multiplyResult_payload_22 = mulOut_22_payload;
  assign io_multiplyResult_payload_23 = mulOut_23_payload;
  assign io_multiplyResult_payload_24 = mulOut_24_payload;
  assign io_multiplyResult_payload_25 = mulOut_25_payload;
  assign io_multiplyResult_payload_26 = mulOut_26_payload;
  assign io_multiplyResult_payload_27 = mulOut_27_payload;
  assign io_multiplyResult_payload_28 = mulOut_28_payload;
  assign io_multiplyResult_payload_29 = mulOut_29_payload;
  assign io_multiplyResult_payload_30 = mulOut_30_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      signalInput_0_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_1_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_2_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_3_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_4_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_5_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_6_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_7_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_8_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_9_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_10_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_11_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_12_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_13_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_14_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_15_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_16_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_17_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_18_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_19_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_20_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_21_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_22_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_23_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_24_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_25_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_26_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_27_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_28_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_29_fork_io_outputs_0_rValid <= 1'b0;
      signalInput_30_fork_io_outputs_0_rValid <= 1'b0;
    end else begin
      if(signalInput_0_fork_io_outputs_0_ready) begin
        signalInput_0_fork_io_outputs_0_rValid <= signalInput_0_fork_io_outputs_0_valid;
      end
      if(signalInput_1_fork_io_outputs_0_ready) begin
        signalInput_1_fork_io_outputs_0_rValid <= signalInput_1_fork_io_outputs_0_valid;
      end
      if(signalInput_2_fork_io_outputs_0_ready) begin
        signalInput_2_fork_io_outputs_0_rValid <= signalInput_2_fork_io_outputs_0_valid;
      end
      if(signalInput_3_fork_io_outputs_0_ready) begin
        signalInput_3_fork_io_outputs_0_rValid <= signalInput_3_fork_io_outputs_0_valid;
      end
      if(signalInput_4_fork_io_outputs_0_ready) begin
        signalInput_4_fork_io_outputs_0_rValid <= signalInput_4_fork_io_outputs_0_valid;
      end
      if(signalInput_5_fork_io_outputs_0_ready) begin
        signalInput_5_fork_io_outputs_0_rValid <= signalInput_5_fork_io_outputs_0_valid;
      end
      if(signalInput_6_fork_io_outputs_0_ready) begin
        signalInput_6_fork_io_outputs_0_rValid <= signalInput_6_fork_io_outputs_0_valid;
      end
      if(signalInput_7_fork_io_outputs_0_ready) begin
        signalInput_7_fork_io_outputs_0_rValid <= signalInput_7_fork_io_outputs_0_valid;
      end
      if(signalInput_8_fork_io_outputs_0_ready) begin
        signalInput_8_fork_io_outputs_0_rValid <= signalInput_8_fork_io_outputs_0_valid;
      end
      if(signalInput_9_fork_io_outputs_0_ready) begin
        signalInput_9_fork_io_outputs_0_rValid <= signalInput_9_fork_io_outputs_0_valid;
      end
      if(signalInput_10_fork_io_outputs_0_ready) begin
        signalInput_10_fork_io_outputs_0_rValid <= signalInput_10_fork_io_outputs_0_valid;
      end
      if(signalInput_11_fork_io_outputs_0_ready) begin
        signalInput_11_fork_io_outputs_0_rValid <= signalInput_11_fork_io_outputs_0_valid;
      end
      if(signalInput_12_fork_io_outputs_0_ready) begin
        signalInput_12_fork_io_outputs_0_rValid <= signalInput_12_fork_io_outputs_0_valid;
      end
      if(signalInput_13_fork_io_outputs_0_ready) begin
        signalInput_13_fork_io_outputs_0_rValid <= signalInput_13_fork_io_outputs_0_valid;
      end
      if(signalInput_14_fork_io_outputs_0_ready) begin
        signalInput_14_fork_io_outputs_0_rValid <= signalInput_14_fork_io_outputs_0_valid;
      end
      if(signalInput_15_fork_io_outputs_0_ready) begin
        signalInput_15_fork_io_outputs_0_rValid <= signalInput_15_fork_io_outputs_0_valid;
      end
      if(signalInput_16_fork_io_outputs_0_ready) begin
        signalInput_16_fork_io_outputs_0_rValid <= signalInput_16_fork_io_outputs_0_valid;
      end
      if(signalInput_17_fork_io_outputs_0_ready) begin
        signalInput_17_fork_io_outputs_0_rValid <= signalInput_17_fork_io_outputs_0_valid;
      end
      if(signalInput_18_fork_io_outputs_0_ready) begin
        signalInput_18_fork_io_outputs_0_rValid <= signalInput_18_fork_io_outputs_0_valid;
      end
      if(signalInput_19_fork_io_outputs_0_ready) begin
        signalInput_19_fork_io_outputs_0_rValid <= signalInput_19_fork_io_outputs_0_valid;
      end
      if(signalInput_20_fork_io_outputs_0_ready) begin
        signalInput_20_fork_io_outputs_0_rValid <= signalInput_20_fork_io_outputs_0_valid;
      end
      if(signalInput_21_fork_io_outputs_0_ready) begin
        signalInput_21_fork_io_outputs_0_rValid <= signalInput_21_fork_io_outputs_0_valid;
      end
      if(signalInput_22_fork_io_outputs_0_ready) begin
        signalInput_22_fork_io_outputs_0_rValid <= signalInput_22_fork_io_outputs_0_valid;
      end
      if(signalInput_23_fork_io_outputs_0_ready) begin
        signalInput_23_fork_io_outputs_0_rValid <= signalInput_23_fork_io_outputs_0_valid;
      end
      if(signalInput_24_fork_io_outputs_0_ready) begin
        signalInput_24_fork_io_outputs_0_rValid <= signalInput_24_fork_io_outputs_0_valid;
      end
      if(signalInput_25_fork_io_outputs_0_ready) begin
        signalInput_25_fork_io_outputs_0_rValid <= signalInput_25_fork_io_outputs_0_valid;
      end
      if(signalInput_26_fork_io_outputs_0_ready) begin
        signalInput_26_fork_io_outputs_0_rValid <= signalInput_26_fork_io_outputs_0_valid;
      end
      if(signalInput_27_fork_io_outputs_0_ready) begin
        signalInput_27_fork_io_outputs_0_rValid <= signalInput_27_fork_io_outputs_0_valid;
      end
      if(signalInput_28_fork_io_outputs_0_ready) begin
        signalInput_28_fork_io_outputs_0_rValid <= signalInput_28_fork_io_outputs_0_valid;
      end
      if(signalInput_29_fork_io_outputs_0_ready) begin
        signalInput_29_fork_io_outputs_0_rValid <= signalInput_29_fork_io_outputs_0_valid;
      end
      if(signalInput_30_fork_io_outputs_0_ready) begin
        signalInput_30_fork_io_outputs_0_rValid <= signalInput_30_fork_io_outputs_0_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(signalInput_0_fork_io_outputs_0_ready) begin
      signalInput_0_fork_io_outputs_0_rData <= signalInput_0_fork_io_outputs_0_payload;
    end
    if(signalInput_1_fork_io_outputs_0_ready) begin
      signalInput_1_fork_io_outputs_0_rData <= signalInput_1_fork_io_outputs_0_payload;
    end
    if(signalInput_2_fork_io_outputs_0_ready) begin
      signalInput_2_fork_io_outputs_0_rData <= signalInput_2_fork_io_outputs_0_payload;
    end
    if(signalInput_3_fork_io_outputs_0_ready) begin
      signalInput_3_fork_io_outputs_0_rData <= signalInput_3_fork_io_outputs_0_payload;
    end
    if(signalInput_4_fork_io_outputs_0_ready) begin
      signalInput_4_fork_io_outputs_0_rData <= signalInput_4_fork_io_outputs_0_payload;
    end
    if(signalInput_5_fork_io_outputs_0_ready) begin
      signalInput_5_fork_io_outputs_0_rData <= signalInput_5_fork_io_outputs_0_payload;
    end
    if(signalInput_6_fork_io_outputs_0_ready) begin
      signalInput_6_fork_io_outputs_0_rData <= signalInput_6_fork_io_outputs_0_payload;
    end
    if(signalInput_7_fork_io_outputs_0_ready) begin
      signalInput_7_fork_io_outputs_0_rData <= signalInput_7_fork_io_outputs_0_payload;
    end
    if(signalInput_8_fork_io_outputs_0_ready) begin
      signalInput_8_fork_io_outputs_0_rData <= signalInput_8_fork_io_outputs_0_payload;
    end
    if(signalInput_9_fork_io_outputs_0_ready) begin
      signalInput_9_fork_io_outputs_0_rData <= signalInput_9_fork_io_outputs_0_payload;
    end
    if(signalInput_10_fork_io_outputs_0_ready) begin
      signalInput_10_fork_io_outputs_0_rData <= signalInput_10_fork_io_outputs_0_payload;
    end
    if(signalInput_11_fork_io_outputs_0_ready) begin
      signalInput_11_fork_io_outputs_0_rData <= signalInput_11_fork_io_outputs_0_payload;
    end
    if(signalInput_12_fork_io_outputs_0_ready) begin
      signalInput_12_fork_io_outputs_0_rData <= signalInput_12_fork_io_outputs_0_payload;
    end
    if(signalInput_13_fork_io_outputs_0_ready) begin
      signalInput_13_fork_io_outputs_0_rData <= signalInput_13_fork_io_outputs_0_payload;
    end
    if(signalInput_14_fork_io_outputs_0_ready) begin
      signalInput_14_fork_io_outputs_0_rData <= signalInput_14_fork_io_outputs_0_payload;
    end
    if(signalInput_15_fork_io_outputs_0_ready) begin
      signalInput_15_fork_io_outputs_0_rData <= signalInput_15_fork_io_outputs_0_payload;
    end
    if(signalInput_16_fork_io_outputs_0_ready) begin
      signalInput_16_fork_io_outputs_0_rData <= signalInput_16_fork_io_outputs_0_payload;
    end
    if(signalInput_17_fork_io_outputs_0_ready) begin
      signalInput_17_fork_io_outputs_0_rData <= signalInput_17_fork_io_outputs_0_payload;
    end
    if(signalInput_18_fork_io_outputs_0_ready) begin
      signalInput_18_fork_io_outputs_0_rData <= signalInput_18_fork_io_outputs_0_payload;
    end
    if(signalInput_19_fork_io_outputs_0_ready) begin
      signalInput_19_fork_io_outputs_0_rData <= signalInput_19_fork_io_outputs_0_payload;
    end
    if(signalInput_20_fork_io_outputs_0_ready) begin
      signalInput_20_fork_io_outputs_0_rData <= signalInput_20_fork_io_outputs_0_payload;
    end
    if(signalInput_21_fork_io_outputs_0_ready) begin
      signalInput_21_fork_io_outputs_0_rData <= signalInput_21_fork_io_outputs_0_payload;
    end
    if(signalInput_22_fork_io_outputs_0_ready) begin
      signalInput_22_fork_io_outputs_0_rData <= signalInput_22_fork_io_outputs_0_payload;
    end
    if(signalInput_23_fork_io_outputs_0_ready) begin
      signalInput_23_fork_io_outputs_0_rData <= signalInput_23_fork_io_outputs_0_payload;
    end
    if(signalInput_24_fork_io_outputs_0_ready) begin
      signalInput_24_fork_io_outputs_0_rData <= signalInput_24_fork_io_outputs_0_payload;
    end
    if(signalInput_25_fork_io_outputs_0_ready) begin
      signalInput_25_fork_io_outputs_0_rData <= signalInput_25_fork_io_outputs_0_payload;
    end
    if(signalInput_26_fork_io_outputs_0_ready) begin
      signalInput_26_fork_io_outputs_0_rData <= signalInput_26_fork_io_outputs_0_payload;
    end
    if(signalInput_27_fork_io_outputs_0_ready) begin
      signalInput_27_fork_io_outputs_0_rData <= signalInput_27_fork_io_outputs_0_payload;
    end
    if(signalInput_28_fork_io_outputs_0_ready) begin
      signalInput_28_fork_io_outputs_0_rData <= signalInput_28_fork_io_outputs_0_payload;
    end
    if(signalInput_29_fork_io_outputs_0_ready) begin
      signalInput_29_fork_io_outputs_0_rData <= signalInput_29_fork_io_outputs_0_payload;
    end
    if(signalInput_30_fork_io_outputs_0_ready) begin
      signalInput_30_fork_io_outputs_0_rData <= signalInput_30_fork_io_outputs_0_payload;
    end
  end


endmodule

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

module StreamFork (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload
);

  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload = io_input_payload;
  assign io_outputs_1_payload = io_input_payload;

endmodule
