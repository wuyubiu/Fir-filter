// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : FirSymmetry



module FirSymmetry (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload,
  output              io_output_valid,
  input               io_output_ready,
  output     [21:0]   io_output_payload,
  input               clk,
  input               reset
);
  reg                 inputAll_0_fork_io_outputs_1_ready;
  reg                 inputAll_1_fork_io_outputs_1_ready;
  reg                 inputAll_2_fork_io_outputs_1_ready;
  reg                 inputAll_3_fork_io_outputs_1_ready;
  reg                 inputAll_4_fork_io_outputs_1_ready;
  reg                 inputAll_5_fork_io_outputs_1_ready;
  reg                 inputAll_6_fork_io_outputs_1_ready;
  reg                 inputAll_7_fork_io_outputs_1_ready;
  reg                 inputAll_8_fork_io_outputs_1_ready;
  reg                 inputAll_9_fork_io_outputs_1_ready;
  reg                 inputAll_10_fork_io_outputs_1_ready;
  reg                 inputAll_11_fork_io_outputs_1_ready;
  reg                 inputAll_12_fork_io_outputs_1_ready;
  reg                 inputAll_13_fork_io_outputs_1_ready;
  reg                 inputAll_14_fork_io_outputs_1_ready;
  reg                 inputAll_15_fork_io_outputs_1_ready;
  reg                 inputAll_16_fork_io_outputs_1_ready;
  reg                 inputAll_17_fork_io_outputs_1_ready;
  reg                 inputAll_18_fork_io_outputs_1_ready;
  reg                 inputAll_19_fork_io_outputs_1_ready;
  reg                 inputAll_20_fork_io_outputs_1_ready;
  reg                 inputAll_21_fork_io_outputs_1_ready;
  reg                 inputAll_22_fork_io_outputs_1_ready;
  reg                 inputAll_23_fork_io_outputs_1_ready;
  reg                 inputAll_24_fork_io_outputs_1_ready;
  reg                 inputAll_25_fork_io_outputs_1_ready;
  reg                 inputAll_26_fork_io_outputs_1_ready;
  reg                 inputAll_27_fork_io_outputs_1_ready;
  reg                 inputAll_28_fork_io_outputs_1_ready;
  reg                 inputAll_29_fork_io_outputs_1_ready;
  reg                 inputAll_30_fork_io_outputs_1_ready;
  reg                 inputAll_31_fork_io_outputs_1_ready;
  reg                 inputAll_32_fork_io_outputs_1_ready;
  reg                 inputAll_33_fork_io_outputs_1_ready;
  reg                 inputAll_34_fork_io_outputs_1_ready;
  reg                 inputAll_35_fork_io_outputs_1_ready;
  reg                 inputAll_36_fork_io_outputs_1_ready;
  reg                 inputAll_37_fork_io_outputs_1_ready;
  reg                 inputAll_38_fork_io_outputs_1_ready;
  reg                 inputAll_39_fork_io_outputs_1_ready;
  reg                 inputAll_40_fork_io_outputs_1_ready;
  reg                 inputAll_41_fork_io_outputs_1_ready;
  reg                 inputAll_42_fork_io_outputs_1_ready;
  reg                 inputAll_43_fork_io_outputs_1_ready;
  reg                 inputAll_44_fork_io_outputs_1_ready;
  reg                 inputAll_45_fork_io_outputs_1_ready;
  reg                 inputAll_46_fork_io_outputs_1_ready;
  reg                 inputAll_47_fork_io_outputs_1_ready;
  reg                 inputAll_48_fork_io_outputs_1_ready;
  reg                 inputAll_49_fork_io_outputs_1_ready;
  reg                 inputAll_50_fork_io_outputs_1_ready;
  reg                 inputAll_51_fork_io_outputs_1_ready;
  reg                 inputAll_52_fork_io_outputs_1_ready;
  reg                 inputAll_53_fork_io_outputs_1_ready;
  reg                 inputAll_54_fork_io_outputs_1_ready;
  reg                 inputAll_55_fork_io_outputs_1_ready;
  reg                 inputAll_56_fork_io_outputs_1_ready;
  reg                 inputAll_57_fork_io_outputs_1_ready;
  reg                 inputAll_58_fork_io_outputs_1_ready;
  reg                 inputAll_59_fork_io_outputs_1_ready;
  reg                 inputAll_60_fork_io_outputs_1_ready;
  reg                 inputAll_61_fork_io_outputs_1_ready;
  reg                 inputAll_62_fork_io_outputs_1_ready;
  reg                 inputAll_63_fork_io_outputs_1_ready;
  reg                 inputAll_64_fork_io_outputs_1_ready;
  reg                 inputAll_65_fork_io_outputs_1_ready;
  reg                 inputAll_66_fork_io_outputs_1_ready;
  reg                 inputAll_67_fork_io_outputs_1_ready;
  reg                 inputAll_68_fork_io_outputs_1_ready;
  reg                 inputAll_69_fork_io_outputs_1_ready;
  reg                 inputAll_70_fork_io_outputs_1_ready;
  reg                 inputAll_71_fork_io_outputs_1_ready;
  reg                 inputAll_72_fork_io_outputs_1_ready;
  reg                 inputAll_73_fork_io_outputs_1_ready;
  reg                 inputAll_74_fork_io_outputs_1_ready;
  reg                 inputAll_75_fork_io_outputs_1_ready;
  reg                 inputAll_76_fork_io_outputs_1_ready;
  reg                 inputAll_77_fork_io_outputs_1_ready;
  reg                 inputAll_78_fork_io_outputs_1_ready;
  reg                 inputAll_79_fork_io_outputs_1_ready;
  reg                 inputAll_80_fork_io_outputs_1_ready;
  reg                 inputAll_81_fork_io_outputs_1_ready;
  reg                 inputAll_82_fork_io_outputs_1_ready;
  reg                 inputAll_83_fork_io_outputs_1_ready;
  reg                 inputAll_84_fork_io_outputs_1_ready;
  reg                 inputAll_85_fork_io_outputs_1_ready;
  reg                 inputAll_86_fork_io_outputs_1_ready;
  reg                 inputAll_87_fork_io_outputs_1_ready;
  reg                 inputAll_88_fork_io_outputs_1_ready;
  reg                 inputAll_89_fork_io_outputs_1_ready;
  reg                 inputAll_90_fork_io_outputs_1_ready;
  reg                 inputAll_91_fork_io_outputs_1_ready;
  reg                 inputAll_92_fork_io_outputs_1_ready;
  reg                 inputAll_93_fork_io_outputs_1_ready;
  reg                 inputAll_94_fork_io_outputs_1_ready;
  reg                 inputAll_95_fork_io_outputs_1_ready;
  reg                 inputAll_96_fork_io_outputs_1_ready;
  reg                 inputAll_97_fork_io_outputs_1_ready;
  reg                 inputAll_98_fork_io_outputs_1_ready;
  reg                 inputAll_99_fork_io_outputs_1_ready;
  reg                 inputAll_100_fork_io_outputs_1_ready;
  reg                 inputAll_101_fork_io_outputs_1_ready;
  reg                 inputAll_102_fork_io_outputs_1_ready;
  reg                 inputAll_103_fork_io_outputs_1_ready;
  reg                 inputAll_104_fork_io_outputs_1_ready;
  reg                 inputAll_105_fork_io_outputs_1_ready;
  reg                 inputAll_106_fork_io_outputs_1_ready;
  reg                 inputAll_107_fork_io_outputs_1_ready;
  reg                 inputAll_108_fork_io_outputs_1_ready;
  reg                 inputAll_109_fork_io_outputs_1_ready;
  reg                 inputAll_110_fork_io_outputs_1_ready;
  reg                 inputAll_111_fork_io_outputs_1_ready;
  reg                 inputAll_112_fork_io_outputs_1_ready;
  reg                 inputAll_113_fork_io_outputs_1_ready;
  reg                 inputAll_114_fork_io_outputs_1_ready;
  reg                 inputAll_115_fork_io_outputs_1_ready;
  reg                 inputAll_116_fork_io_outputs_1_ready;
  reg                 inputAll_117_fork_io_outputs_1_ready;
  reg                 inputAll_118_fork_io_outputs_1_ready;
  reg                 inputAll_119_fork_io_outputs_1_ready;
  reg                 inputAll_120_fork_io_outputs_1_ready;
  reg                 inputAll_121_fork_io_outputs_1_ready;
  reg                 inputAll_122_fork_io_outputs_1_ready;
  reg                 inputAll_123_fork_io_outputs_1_ready;
  reg                 inputAll_124_fork_io_outputs_1_ready;
  reg                 inputAll_125_fork_io_outputs_1_ready;
  reg                 inputAll_126_fork_io_outputs_1_ready;
  reg                 inputAll_127_fork_io_outputs_1_ready;
  wire                inputAll_0_fork_io_input_ready;
  wire                inputAll_0_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_0_fork_io_outputs_0_payload;
  wire                inputAll_0_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_0_fork_io_outputs_1_payload;
  wire                inputAll_1_fork_io_input_ready;
  wire                inputAll_1_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_1_fork_io_outputs_0_payload;
  wire                inputAll_1_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_1_fork_io_outputs_1_payload;
  wire                inputAll_2_fork_io_input_ready;
  wire                inputAll_2_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_2_fork_io_outputs_0_payload;
  wire                inputAll_2_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_2_fork_io_outputs_1_payload;
  wire                inputAll_3_fork_io_input_ready;
  wire                inputAll_3_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_3_fork_io_outputs_0_payload;
  wire                inputAll_3_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_3_fork_io_outputs_1_payload;
  wire                inputAll_4_fork_io_input_ready;
  wire                inputAll_4_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_4_fork_io_outputs_0_payload;
  wire                inputAll_4_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_4_fork_io_outputs_1_payload;
  wire                inputAll_5_fork_io_input_ready;
  wire                inputAll_5_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_5_fork_io_outputs_0_payload;
  wire                inputAll_5_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_5_fork_io_outputs_1_payload;
  wire                inputAll_6_fork_io_input_ready;
  wire                inputAll_6_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_6_fork_io_outputs_0_payload;
  wire                inputAll_6_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_6_fork_io_outputs_1_payload;
  wire                inputAll_7_fork_io_input_ready;
  wire                inputAll_7_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_7_fork_io_outputs_0_payload;
  wire                inputAll_7_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_7_fork_io_outputs_1_payload;
  wire                inputAll_8_fork_io_input_ready;
  wire                inputAll_8_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_8_fork_io_outputs_0_payload;
  wire                inputAll_8_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_8_fork_io_outputs_1_payload;
  wire                inputAll_9_fork_io_input_ready;
  wire                inputAll_9_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_9_fork_io_outputs_0_payload;
  wire                inputAll_9_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_9_fork_io_outputs_1_payload;
  wire                inputAll_10_fork_io_input_ready;
  wire                inputAll_10_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_10_fork_io_outputs_0_payload;
  wire                inputAll_10_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_10_fork_io_outputs_1_payload;
  wire                inputAll_11_fork_io_input_ready;
  wire                inputAll_11_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_11_fork_io_outputs_0_payload;
  wire                inputAll_11_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_11_fork_io_outputs_1_payload;
  wire                inputAll_12_fork_io_input_ready;
  wire                inputAll_12_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_12_fork_io_outputs_0_payload;
  wire                inputAll_12_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_12_fork_io_outputs_1_payload;
  wire                inputAll_13_fork_io_input_ready;
  wire                inputAll_13_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_13_fork_io_outputs_0_payload;
  wire                inputAll_13_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_13_fork_io_outputs_1_payload;
  wire                inputAll_14_fork_io_input_ready;
  wire                inputAll_14_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_14_fork_io_outputs_0_payload;
  wire                inputAll_14_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_14_fork_io_outputs_1_payload;
  wire                inputAll_15_fork_io_input_ready;
  wire                inputAll_15_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_15_fork_io_outputs_0_payload;
  wire                inputAll_15_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_15_fork_io_outputs_1_payload;
  wire                inputAll_16_fork_io_input_ready;
  wire                inputAll_16_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_16_fork_io_outputs_0_payload;
  wire                inputAll_16_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_16_fork_io_outputs_1_payload;
  wire                inputAll_17_fork_io_input_ready;
  wire                inputAll_17_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_17_fork_io_outputs_0_payload;
  wire                inputAll_17_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_17_fork_io_outputs_1_payload;
  wire                inputAll_18_fork_io_input_ready;
  wire                inputAll_18_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_18_fork_io_outputs_0_payload;
  wire                inputAll_18_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_18_fork_io_outputs_1_payload;
  wire                inputAll_19_fork_io_input_ready;
  wire                inputAll_19_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_19_fork_io_outputs_0_payload;
  wire                inputAll_19_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_19_fork_io_outputs_1_payload;
  wire                inputAll_20_fork_io_input_ready;
  wire                inputAll_20_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_20_fork_io_outputs_0_payload;
  wire                inputAll_20_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_20_fork_io_outputs_1_payload;
  wire                inputAll_21_fork_io_input_ready;
  wire                inputAll_21_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_21_fork_io_outputs_0_payload;
  wire                inputAll_21_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_21_fork_io_outputs_1_payload;
  wire                inputAll_22_fork_io_input_ready;
  wire                inputAll_22_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_22_fork_io_outputs_0_payload;
  wire                inputAll_22_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_22_fork_io_outputs_1_payload;
  wire                inputAll_23_fork_io_input_ready;
  wire                inputAll_23_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_23_fork_io_outputs_0_payload;
  wire                inputAll_23_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_23_fork_io_outputs_1_payload;
  wire                inputAll_24_fork_io_input_ready;
  wire                inputAll_24_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_24_fork_io_outputs_0_payload;
  wire                inputAll_24_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_24_fork_io_outputs_1_payload;
  wire                inputAll_25_fork_io_input_ready;
  wire                inputAll_25_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_25_fork_io_outputs_0_payload;
  wire                inputAll_25_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_25_fork_io_outputs_1_payload;
  wire                inputAll_26_fork_io_input_ready;
  wire                inputAll_26_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_26_fork_io_outputs_0_payload;
  wire                inputAll_26_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_26_fork_io_outputs_1_payload;
  wire                inputAll_27_fork_io_input_ready;
  wire                inputAll_27_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_27_fork_io_outputs_0_payload;
  wire                inputAll_27_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_27_fork_io_outputs_1_payload;
  wire                inputAll_28_fork_io_input_ready;
  wire                inputAll_28_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_28_fork_io_outputs_0_payload;
  wire                inputAll_28_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_28_fork_io_outputs_1_payload;
  wire                inputAll_29_fork_io_input_ready;
  wire                inputAll_29_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_29_fork_io_outputs_0_payload;
  wire                inputAll_29_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_29_fork_io_outputs_1_payload;
  wire                inputAll_30_fork_io_input_ready;
  wire                inputAll_30_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_30_fork_io_outputs_0_payload;
  wire                inputAll_30_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_30_fork_io_outputs_1_payload;
  wire                inputAll_31_fork_io_input_ready;
  wire                inputAll_31_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_31_fork_io_outputs_0_payload;
  wire                inputAll_31_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_31_fork_io_outputs_1_payload;
  wire                inputAll_32_fork_io_input_ready;
  wire                inputAll_32_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_32_fork_io_outputs_0_payload;
  wire                inputAll_32_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_32_fork_io_outputs_1_payload;
  wire                inputAll_33_fork_io_input_ready;
  wire                inputAll_33_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_33_fork_io_outputs_0_payload;
  wire                inputAll_33_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_33_fork_io_outputs_1_payload;
  wire                inputAll_34_fork_io_input_ready;
  wire                inputAll_34_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_34_fork_io_outputs_0_payload;
  wire                inputAll_34_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_34_fork_io_outputs_1_payload;
  wire                inputAll_35_fork_io_input_ready;
  wire                inputAll_35_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_35_fork_io_outputs_0_payload;
  wire                inputAll_35_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_35_fork_io_outputs_1_payload;
  wire                inputAll_36_fork_io_input_ready;
  wire                inputAll_36_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_36_fork_io_outputs_0_payload;
  wire                inputAll_36_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_36_fork_io_outputs_1_payload;
  wire                inputAll_37_fork_io_input_ready;
  wire                inputAll_37_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_37_fork_io_outputs_0_payload;
  wire                inputAll_37_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_37_fork_io_outputs_1_payload;
  wire                inputAll_38_fork_io_input_ready;
  wire                inputAll_38_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_38_fork_io_outputs_0_payload;
  wire                inputAll_38_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_38_fork_io_outputs_1_payload;
  wire                inputAll_39_fork_io_input_ready;
  wire                inputAll_39_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_39_fork_io_outputs_0_payload;
  wire                inputAll_39_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_39_fork_io_outputs_1_payload;
  wire                inputAll_40_fork_io_input_ready;
  wire                inputAll_40_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_40_fork_io_outputs_0_payload;
  wire                inputAll_40_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_40_fork_io_outputs_1_payload;
  wire                inputAll_41_fork_io_input_ready;
  wire                inputAll_41_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_41_fork_io_outputs_0_payload;
  wire                inputAll_41_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_41_fork_io_outputs_1_payload;
  wire                inputAll_42_fork_io_input_ready;
  wire                inputAll_42_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_42_fork_io_outputs_0_payload;
  wire                inputAll_42_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_42_fork_io_outputs_1_payload;
  wire                inputAll_43_fork_io_input_ready;
  wire                inputAll_43_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_43_fork_io_outputs_0_payload;
  wire                inputAll_43_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_43_fork_io_outputs_1_payload;
  wire                inputAll_44_fork_io_input_ready;
  wire                inputAll_44_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_44_fork_io_outputs_0_payload;
  wire                inputAll_44_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_44_fork_io_outputs_1_payload;
  wire                inputAll_45_fork_io_input_ready;
  wire                inputAll_45_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_45_fork_io_outputs_0_payload;
  wire                inputAll_45_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_45_fork_io_outputs_1_payload;
  wire                inputAll_46_fork_io_input_ready;
  wire                inputAll_46_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_46_fork_io_outputs_0_payload;
  wire                inputAll_46_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_46_fork_io_outputs_1_payload;
  wire                inputAll_47_fork_io_input_ready;
  wire                inputAll_47_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_47_fork_io_outputs_0_payload;
  wire                inputAll_47_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_47_fork_io_outputs_1_payload;
  wire                inputAll_48_fork_io_input_ready;
  wire                inputAll_48_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_48_fork_io_outputs_0_payload;
  wire                inputAll_48_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_48_fork_io_outputs_1_payload;
  wire                inputAll_49_fork_io_input_ready;
  wire                inputAll_49_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_49_fork_io_outputs_0_payload;
  wire                inputAll_49_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_49_fork_io_outputs_1_payload;
  wire                inputAll_50_fork_io_input_ready;
  wire                inputAll_50_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_50_fork_io_outputs_0_payload;
  wire                inputAll_50_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_50_fork_io_outputs_1_payload;
  wire                inputAll_51_fork_io_input_ready;
  wire                inputAll_51_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_51_fork_io_outputs_0_payload;
  wire                inputAll_51_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_51_fork_io_outputs_1_payload;
  wire                inputAll_52_fork_io_input_ready;
  wire                inputAll_52_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_52_fork_io_outputs_0_payload;
  wire                inputAll_52_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_52_fork_io_outputs_1_payload;
  wire                inputAll_53_fork_io_input_ready;
  wire                inputAll_53_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_53_fork_io_outputs_0_payload;
  wire                inputAll_53_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_53_fork_io_outputs_1_payload;
  wire                inputAll_54_fork_io_input_ready;
  wire                inputAll_54_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_54_fork_io_outputs_0_payload;
  wire                inputAll_54_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_54_fork_io_outputs_1_payload;
  wire                inputAll_55_fork_io_input_ready;
  wire                inputAll_55_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_55_fork_io_outputs_0_payload;
  wire                inputAll_55_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_55_fork_io_outputs_1_payload;
  wire                inputAll_56_fork_io_input_ready;
  wire                inputAll_56_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_56_fork_io_outputs_0_payload;
  wire                inputAll_56_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_56_fork_io_outputs_1_payload;
  wire                inputAll_57_fork_io_input_ready;
  wire                inputAll_57_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_57_fork_io_outputs_0_payload;
  wire                inputAll_57_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_57_fork_io_outputs_1_payload;
  wire                inputAll_58_fork_io_input_ready;
  wire                inputAll_58_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_58_fork_io_outputs_0_payload;
  wire                inputAll_58_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_58_fork_io_outputs_1_payload;
  wire                inputAll_59_fork_io_input_ready;
  wire                inputAll_59_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_59_fork_io_outputs_0_payload;
  wire                inputAll_59_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_59_fork_io_outputs_1_payload;
  wire                inputAll_60_fork_io_input_ready;
  wire                inputAll_60_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_60_fork_io_outputs_0_payload;
  wire                inputAll_60_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_60_fork_io_outputs_1_payload;
  wire                inputAll_61_fork_io_input_ready;
  wire                inputAll_61_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_61_fork_io_outputs_0_payload;
  wire                inputAll_61_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_61_fork_io_outputs_1_payload;
  wire                inputAll_62_fork_io_input_ready;
  wire                inputAll_62_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_62_fork_io_outputs_0_payload;
  wire                inputAll_62_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_62_fork_io_outputs_1_payload;
  wire                inputAll_63_fork_io_input_ready;
  wire                inputAll_63_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_63_fork_io_outputs_0_payload;
  wire                inputAll_63_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_63_fork_io_outputs_1_payload;
  wire                inputAll_64_fork_io_input_ready;
  wire                inputAll_64_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_64_fork_io_outputs_0_payload;
  wire                inputAll_64_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_64_fork_io_outputs_1_payload;
  wire                inputAll_65_fork_io_input_ready;
  wire                inputAll_65_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_65_fork_io_outputs_0_payload;
  wire                inputAll_65_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_65_fork_io_outputs_1_payload;
  wire                inputAll_66_fork_io_input_ready;
  wire                inputAll_66_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_66_fork_io_outputs_0_payload;
  wire                inputAll_66_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_66_fork_io_outputs_1_payload;
  wire                inputAll_67_fork_io_input_ready;
  wire                inputAll_67_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_67_fork_io_outputs_0_payload;
  wire                inputAll_67_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_67_fork_io_outputs_1_payload;
  wire                inputAll_68_fork_io_input_ready;
  wire                inputAll_68_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_68_fork_io_outputs_0_payload;
  wire                inputAll_68_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_68_fork_io_outputs_1_payload;
  wire                inputAll_69_fork_io_input_ready;
  wire                inputAll_69_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_69_fork_io_outputs_0_payload;
  wire                inputAll_69_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_69_fork_io_outputs_1_payload;
  wire                inputAll_70_fork_io_input_ready;
  wire                inputAll_70_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_70_fork_io_outputs_0_payload;
  wire                inputAll_70_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_70_fork_io_outputs_1_payload;
  wire                inputAll_71_fork_io_input_ready;
  wire                inputAll_71_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_71_fork_io_outputs_0_payload;
  wire                inputAll_71_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_71_fork_io_outputs_1_payload;
  wire                inputAll_72_fork_io_input_ready;
  wire                inputAll_72_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_72_fork_io_outputs_0_payload;
  wire                inputAll_72_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_72_fork_io_outputs_1_payload;
  wire                inputAll_73_fork_io_input_ready;
  wire                inputAll_73_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_73_fork_io_outputs_0_payload;
  wire                inputAll_73_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_73_fork_io_outputs_1_payload;
  wire                inputAll_74_fork_io_input_ready;
  wire                inputAll_74_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_74_fork_io_outputs_0_payload;
  wire                inputAll_74_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_74_fork_io_outputs_1_payload;
  wire                inputAll_75_fork_io_input_ready;
  wire                inputAll_75_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_75_fork_io_outputs_0_payload;
  wire                inputAll_75_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_75_fork_io_outputs_1_payload;
  wire                inputAll_76_fork_io_input_ready;
  wire                inputAll_76_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_76_fork_io_outputs_0_payload;
  wire                inputAll_76_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_76_fork_io_outputs_1_payload;
  wire                inputAll_77_fork_io_input_ready;
  wire                inputAll_77_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_77_fork_io_outputs_0_payload;
  wire                inputAll_77_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_77_fork_io_outputs_1_payload;
  wire                inputAll_78_fork_io_input_ready;
  wire                inputAll_78_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_78_fork_io_outputs_0_payload;
  wire                inputAll_78_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_78_fork_io_outputs_1_payload;
  wire                inputAll_79_fork_io_input_ready;
  wire                inputAll_79_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_79_fork_io_outputs_0_payload;
  wire                inputAll_79_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_79_fork_io_outputs_1_payload;
  wire                inputAll_80_fork_io_input_ready;
  wire                inputAll_80_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_80_fork_io_outputs_0_payload;
  wire                inputAll_80_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_80_fork_io_outputs_1_payload;
  wire                inputAll_81_fork_io_input_ready;
  wire                inputAll_81_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_81_fork_io_outputs_0_payload;
  wire                inputAll_81_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_81_fork_io_outputs_1_payload;
  wire                inputAll_82_fork_io_input_ready;
  wire                inputAll_82_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_82_fork_io_outputs_0_payload;
  wire                inputAll_82_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_82_fork_io_outputs_1_payload;
  wire                inputAll_83_fork_io_input_ready;
  wire                inputAll_83_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_83_fork_io_outputs_0_payload;
  wire                inputAll_83_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_83_fork_io_outputs_1_payload;
  wire                inputAll_84_fork_io_input_ready;
  wire                inputAll_84_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_84_fork_io_outputs_0_payload;
  wire                inputAll_84_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_84_fork_io_outputs_1_payload;
  wire                inputAll_85_fork_io_input_ready;
  wire                inputAll_85_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_85_fork_io_outputs_0_payload;
  wire                inputAll_85_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_85_fork_io_outputs_1_payload;
  wire                inputAll_86_fork_io_input_ready;
  wire                inputAll_86_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_86_fork_io_outputs_0_payload;
  wire                inputAll_86_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_86_fork_io_outputs_1_payload;
  wire                inputAll_87_fork_io_input_ready;
  wire                inputAll_87_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_87_fork_io_outputs_0_payload;
  wire                inputAll_87_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_87_fork_io_outputs_1_payload;
  wire                inputAll_88_fork_io_input_ready;
  wire                inputAll_88_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_88_fork_io_outputs_0_payload;
  wire                inputAll_88_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_88_fork_io_outputs_1_payload;
  wire                inputAll_89_fork_io_input_ready;
  wire                inputAll_89_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_89_fork_io_outputs_0_payload;
  wire                inputAll_89_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_89_fork_io_outputs_1_payload;
  wire                inputAll_90_fork_io_input_ready;
  wire                inputAll_90_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_90_fork_io_outputs_0_payload;
  wire                inputAll_90_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_90_fork_io_outputs_1_payload;
  wire                inputAll_91_fork_io_input_ready;
  wire                inputAll_91_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_91_fork_io_outputs_0_payload;
  wire                inputAll_91_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_91_fork_io_outputs_1_payload;
  wire                inputAll_92_fork_io_input_ready;
  wire                inputAll_92_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_92_fork_io_outputs_0_payload;
  wire                inputAll_92_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_92_fork_io_outputs_1_payload;
  wire                inputAll_93_fork_io_input_ready;
  wire                inputAll_93_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_93_fork_io_outputs_0_payload;
  wire                inputAll_93_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_93_fork_io_outputs_1_payload;
  wire                inputAll_94_fork_io_input_ready;
  wire                inputAll_94_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_94_fork_io_outputs_0_payload;
  wire                inputAll_94_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_94_fork_io_outputs_1_payload;
  wire                inputAll_95_fork_io_input_ready;
  wire                inputAll_95_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_95_fork_io_outputs_0_payload;
  wire                inputAll_95_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_95_fork_io_outputs_1_payload;
  wire                inputAll_96_fork_io_input_ready;
  wire                inputAll_96_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_96_fork_io_outputs_0_payload;
  wire                inputAll_96_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_96_fork_io_outputs_1_payload;
  wire                inputAll_97_fork_io_input_ready;
  wire                inputAll_97_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_97_fork_io_outputs_0_payload;
  wire                inputAll_97_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_97_fork_io_outputs_1_payload;
  wire                inputAll_98_fork_io_input_ready;
  wire                inputAll_98_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_98_fork_io_outputs_0_payload;
  wire                inputAll_98_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_98_fork_io_outputs_1_payload;
  wire                inputAll_99_fork_io_input_ready;
  wire                inputAll_99_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_99_fork_io_outputs_0_payload;
  wire                inputAll_99_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_99_fork_io_outputs_1_payload;
  wire                inputAll_100_fork_io_input_ready;
  wire                inputAll_100_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_100_fork_io_outputs_0_payload;
  wire                inputAll_100_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_100_fork_io_outputs_1_payload;
  wire                inputAll_101_fork_io_input_ready;
  wire                inputAll_101_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_101_fork_io_outputs_0_payload;
  wire                inputAll_101_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_101_fork_io_outputs_1_payload;
  wire                inputAll_102_fork_io_input_ready;
  wire                inputAll_102_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_102_fork_io_outputs_0_payload;
  wire                inputAll_102_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_102_fork_io_outputs_1_payload;
  wire                inputAll_103_fork_io_input_ready;
  wire                inputAll_103_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_103_fork_io_outputs_0_payload;
  wire                inputAll_103_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_103_fork_io_outputs_1_payload;
  wire                inputAll_104_fork_io_input_ready;
  wire                inputAll_104_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_104_fork_io_outputs_0_payload;
  wire                inputAll_104_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_104_fork_io_outputs_1_payload;
  wire                inputAll_105_fork_io_input_ready;
  wire                inputAll_105_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_105_fork_io_outputs_0_payload;
  wire                inputAll_105_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_105_fork_io_outputs_1_payload;
  wire                inputAll_106_fork_io_input_ready;
  wire                inputAll_106_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_106_fork_io_outputs_0_payload;
  wire                inputAll_106_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_106_fork_io_outputs_1_payload;
  wire                inputAll_107_fork_io_input_ready;
  wire                inputAll_107_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_107_fork_io_outputs_0_payload;
  wire                inputAll_107_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_107_fork_io_outputs_1_payload;
  wire                inputAll_108_fork_io_input_ready;
  wire                inputAll_108_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_108_fork_io_outputs_0_payload;
  wire                inputAll_108_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_108_fork_io_outputs_1_payload;
  wire                inputAll_109_fork_io_input_ready;
  wire                inputAll_109_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_109_fork_io_outputs_0_payload;
  wire                inputAll_109_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_109_fork_io_outputs_1_payload;
  wire                inputAll_110_fork_io_input_ready;
  wire                inputAll_110_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_110_fork_io_outputs_0_payload;
  wire                inputAll_110_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_110_fork_io_outputs_1_payload;
  wire                inputAll_111_fork_io_input_ready;
  wire                inputAll_111_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_111_fork_io_outputs_0_payload;
  wire                inputAll_111_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_111_fork_io_outputs_1_payload;
  wire                inputAll_112_fork_io_input_ready;
  wire                inputAll_112_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_112_fork_io_outputs_0_payload;
  wire                inputAll_112_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_112_fork_io_outputs_1_payload;
  wire                inputAll_113_fork_io_input_ready;
  wire                inputAll_113_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_113_fork_io_outputs_0_payload;
  wire                inputAll_113_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_113_fork_io_outputs_1_payload;
  wire                inputAll_114_fork_io_input_ready;
  wire                inputAll_114_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_114_fork_io_outputs_0_payload;
  wire                inputAll_114_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_114_fork_io_outputs_1_payload;
  wire                inputAll_115_fork_io_input_ready;
  wire                inputAll_115_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_115_fork_io_outputs_0_payload;
  wire                inputAll_115_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_115_fork_io_outputs_1_payload;
  wire                inputAll_116_fork_io_input_ready;
  wire                inputAll_116_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_116_fork_io_outputs_0_payload;
  wire                inputAll_116_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_116_fork_io_outputs_1_payload;
  wire                inputAll_117_fork_io_input_ready;
  wire                inputAll_117_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_117_fork_io_outputs_0_payload;
  wire                inputAll_117_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_117_fork_io_outputs_1_payload;
  wire                inputAll_118_fork_io_input_ready;
  wire                inputAll_118_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_118_fork_io_outputs_0_payload;
  wire                inputAll_118_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_118_fork_io_outputs_1_payload;
  wire                inputAll_119_fork_io_input_ready;
  wire                inputAll_119_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_119_fork_io_outputs_0_payload;
  wire                inputAll_119_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_119_fork_io_outputs_1_payload;
  wire                inputAll_120_fork_io_input_ready;
  wire                inputAll_120_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_120_fork_io_outputs_0_payload;
  wire                inputAll_120_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_120_fork_io_outputs_1_payload;
  wire                inputAll_121_fork_io_input_ready;
  wire                inputAll_121_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_121_fork_io_outputs_0_payload;
  wire                inputAll_121_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_121_fork_io_outputs_1_payload;
  wire                inputAll_122_fork_io_input_ready;
  wire                inputAll_122_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_122_fork_io_outputs_0_payload;
  wire                inputAll_122_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_122_fork_io_outputs_1_payload;
  wire                inputAll_123_fork_io_input_ready;
  wire                inputAll_123_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_123_fork_io_outputs_0_payload;
  wire                inputAll_123_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_123_fork_io_outputs_1_payload;
  wire                inputAll_124_fork_io_input_ready;
  wire                inputAll_124_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_124_fork_io_outputs_0_payload;
  wire                inputAll_124_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_124_fork_io_outputs_1_payload;
  wire                inputAll_125_fork_io_input_ready;
  wire                inputAll_125_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_125_fork_io_outputs_0_payload;
  wire                inputAll_125_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_125_fork_io_outputs_1_payload;
  wire                inputAll_126_fork_io_input_ready;
  wire                inputAll_126_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_126_fork_io_outputs_0_payload;
  wire                inputAll_126_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_126_fork_io_outputs_1_payload;
  wire                inputAll_127_fork_io_input_ready;
  wire                inputAll_127_fork_io_outputs_0_valid;
  wire       [7:0]    inputAll_127_fork_io_outputs_0_payload;
  wire                inputAll_127_fork_io_outputs_1_valid;
  wire       [7:0]    inputAll_127_fork_io_outputs_1_payload;
  wire       [8:0]    _zz_mulResGroup_0_payload;
  wire       [8:0]    _zz_mulResGroup_1_payload;
  wire       [8:0]    _zz_mulResGroup_2_payload;
  wire       [8:0]    _zz_mulResGroup_3_payload;
  wire       [8:0]    _zz_mulResGroup_4_payload;
  wire       [8:0]    _zz_mulResGroup_5_payload;
  wire       [8:0]    _zz_mulResGroup_6_payload;
  wire       [8:0]    _zz_mulResGroup_7_payload;
  wire       [8:0]    _zz_mulResGroup_8_payload;
  wire       [8:0]    _zz_mulResGroup_9_payload;
  wire       [8:0]    _zz_mulResGroup_10_payload;
  wire       [8:0]    _zz_mulResGroup_11_payload;
  wire       [8:0]    _zz_mulResGroup_12_payload;
  wire       [8:0]    _zz_mulResGroup_13_payload;
  wire       [8:0]    _zz_mulResGroup_14_payload;
  wire       [8:0]    _zz_mulResGroup_15_payload;
  wire       [9:0]    _zz_mulResGroup_16_payload;
  wire       [0:0]    _zz_mulResGroup_16_payload_1;
  wire       [8:0]    _zz_mulResGroup_16_payload_2;
  wire       [8:0]    _zz_mulResGroup_16_payload_3;
  wire       [8:0]    _zz_mulResGroup_16_payload_4;
  wire       [9:0]    _zz_mulResGroup_17_payload;
  wire       [0:0]    _zz_mulResGroup_17_payload_1;
  wire       [8:0]    _zz_mulResGroup_17_payload_2;
  wire       [8:0]    _zz_mulResGroup_17_payload_3;
  wire       [8:0]    _zz_mulResGroup_17_payload_4;
  wire       [9:0]    _zz_mulResGroup_18_payload;
  wire       [0:0]    _zz_mulResGroup_18_payload_1;
  wire       [8:0]    _zz_mulResGroup_18_payload_2;
  wire       [8:0]    _zz_mulResGroup_18_payload_3;
  wire       [8:0]    _zz_mulResGroup_18_payload_4;
  wire       [8:0]    _zz_mulResGroup_19_payload;
  wire       [8:0]    _zz_mulResGroup_20_payload;
  wire       [10:0]   _zz_mulResGroup_21_payload;
  wire       [1:0]    _zz_mulResGroup_21_payload_1;
  wire       [8:0]    _zz_mulResGroup_21_payload_2;
  wire       [8:0]    _zz_mulResGroup_21_payload_3;
  wire       [8:0]    _zz_mulResGroup_21_payload_4;
  wire       [10:0]   _zz_mulResGroup_22_payload;
  wire       [1:0]    _zz_mulResGroup_22_payload_1;
  wire       [8:0]    _zz_mulResGroup_22_payload_2;
  wire       [8:0]    _zz_mulResGroup_22_payload_3;
  wire       [8:0]    _zz_mulResGroup_22_payload_4;
  wire       [10:0]   _zz_mulResGroup_23_payload;
  wire       [1:0]    _zz_mulResGroup_23_payload_1;
  wire       [8:0]    _zz_mulResGroup_23_payload_2;
  wire       [8:0]    _zz_mulResGroup_23_payload_3;
  wire       [8:0]    _zz_mulResGroup_23_payload_4;
  wire       [10:0]   _zz_mulResGroup_24_payload;
  wire       [1:0]    _zz_mulResGroup_24_payload_1;
  wire       [8:0]    _zz_mulResGroup_24_payload_2;
  wire       [8:0]    _zz_mulResGroup_24_payload_3;
  wire       [8:0]    _zz_mulResGroup_24_payload_4;
  wire       [10:0]   _zz_mulResGroup_25_payload;
  wire       [1:0]    _zz_mulResGroup_25_payload_1;
  wire       [8:0]    _zz_mulResGroup_25_payload_2;
  wire       [8:0]    _zz_mulResGroup_25_payload_3;
  wire       [8:0]    _zz_mulResGroup_25_payload_4;
  wire       [8:0]    _zz_mulResGroup_26_payload;
  wire       [9:0]    _zz_mulResGroup_27_payload;
  wire       [0:0]    _zz_mulResGroup_27_payload_1;
  wire       [8:0]    _zz_mulResGroup_27_payload_2;
  wire       [8:0]    _zz_mulResGroup_27_payload_3;
  wire       [8:0]    _zz_mulResGroup_27_payload_4;
  wire       [10:0]   _zz_mulResGroup_28_payload;
  wire       [1:0]    _zz_mulResGroup_28_payload_1;
  wire       [8:0]    _zz_mulResGroup_28_payload_2;
  wire       [8:0]    _zz_mulResGroup_28_payload_3;
  wire       [8:0]    _zz_mulResGroup_28_payload_4;
  wire       [10:0]   _zz_mulResGroup_29_payload;
  wire       [1:0]    _zz_mulResGroup_29_payload_1;
  wire       [8:0]    _zz_mulResGroup_29_payload_2;
  wire       [8:0]    _zz_mulResGroup_29_payload_3;
  wire       [8:0]    _zz_mulResGroup_29_payload_4;
  wire       [10:0]   _zz_mulResGroup_30_payload;
  wire       [1:0]    _zz_mulResGroup_30_payload_1;
  wire       [8:0]    _zz_mulResGroup_30_payload_2;
  wire       [8:0]    _zz_mulResGroup_30_payload_3;
  wire       [8:0]    _zz_mulResGroup_30_payload_4;
  wire       [10:0]   _zz_mulResGroup_31_payload;
  wire       [1:0]    _zz_mulResGroup_31_payload_1;
  wire       [8:0]    _zz_mulResGroup_31_payload_2;
  wire       [8:0]    _zz_mulResGroup_31_payload_3;
  wire       [8:0]    _zz_mulResGroup_31_payload_4;
  wire       [8:0]    _zz_mulResGroup_32_payload;
  wire       [10:0]   _zz_mulResGroup_33_payload;
  wire       [1:0]    _zz_mulResGroup_33_payload_1;
  wire       [8:0]    _zz_mulResGroup_33_payload_2;
  wire       [8:0]    _zz_mulResGroup_33_payload_3;
  wire       [8:0]    _zz_mulResGroup_33_payload_4;
  wire       [11:0]   _zz_mulResGroup_34_payload;
  wire       [2:0]    _zz_mulResGroup_34_payload_1;
  wire       [8:0]    _zz_mulResGroup_34_payload_2;
  wire       [8:0]    _zz_mulResGroup_34_payload_3;
  wire       [8:0]    _zz_mulResGroup_34_payload_4;
  wire       [11:0]   _zz_mulResGroup_35_payload;
  wire       [2:0]    _zz_mulResGroup_35_payload_1;
  wire       [8:0]    _zz_mulResGroup_35_payload_2;
  wire       [8:0]    _zz_mulResGroup_35_payload_3;
  wire       [8:0]    _zz_mulResGroup_35_payload_4;
  wire       [12:0]   _zz_mulResGroup_36_payload;
  wire       [3:0]    _zz_mulResGroup_36_payload_1;
  wire       [8:0]    _zz_mulResGroup_36_payload_2;
  wire       [8:0]    _zz_mulResGroup_36_payload_3;
  wire       [8:0]    _zz_mulResGroup_36_payload_4;
  wire       [11:0]   _zz_mulResGroup_37_payload;
  wire       [2:0]    _zz_mulResGroup_37_payload_1;
  wire       [8:0]    _zz_mulResGroup_37_payload_2;
  wire       [8:0]    _zz_mulResGroup_37_payload_3;
  wire       [8:0]    _zz_mulResGroup_37_payload_4;
  wire       [10:0]   _zz_mulResGroup_38_payload;
  wire       [1:0]    _zz_mulResGroup_38_payload_1;
  wire       [8:0]    _zz_mulResGroup_38_payload_2;
  wire       [8:0]    _zz_mulResGroup_38_payload_3;
  wire       [8:0]    _zz_mulResGroup_38_payload_4;
  wire       [9:0]    _zz_mulResGroup_39_payload;
  wire       [0:0]    _zz_mulResGroup_39_payload_1;
  wire       [8:0]    _zz_mulResGroup_39_payload_2;
  wire       [8:0]    _zz_mulResGroup_39_payload_3;
  wire       [8:0]    _zz_mulResGroup_39_payload_4;
  wire       [11:0]   _zz_mulResGroup_40_payload;
  wire       [2:0]    _zz_mulResGroup_40_payload_1;
  wire       [8:0]    _zz_mulResGroup_40_payload_2;
  wire       [8:0]    _zz_mulResGroup_40_payload_3;
  wire       [8:0]    _zz_mulResGroup_40_payload_4;
  wire       [12:0]   _zz_mulResGroup_41_payload;
  wire       [3:0]    _zz_mulResGroup_41_payload_1;
  wire       [8:0]    _zz_mulResGroup_41_payload_2;
  wire       [8:0]    _zz_mulResGroup_41_payload_3;
  wire       [8:0]    _zz_mulResGroup_41_payload_4;
  wire       [12:0]   _zz_mulResGroup_42_payload;
  wire       [3:0]    _zz_mulResGroup_42_payload_1;
  wire       [8:0]    _zz_mulResGroup_42_payload_2;
  wire       [8:0]    _zz_mulResGroup_42_payload_3;
  wire       [8:0]    _zz_mulResGroup_42_payload_4;
  wire       [12:0]   _zz_mulResGroup_43_payload;
  wire       [3:0]    _zz_mulResGroup_43_payload_1;
  wire       [8:0]    _zz_mulResGroup_43_payload_2;
  wire       [8:0]    _zz_mulResGroup_43_payload_3;
  wire       [8:0]    _zz_mulResGroup_43_payload_4;
  wire       [10:0]   _zz_mulResGroup_44_payload;
  wire       [1:0]    _zz_mulResGroup_44_payload_1;
  wire       [8:0]    _zz_mulResGroup_44_payload_2;
  wire       [8:0]    _zz_mulResGroup_44_payload_3;
  wire       [8:0]    _zz_mulResGroup_44_payload_4;
  wire       [10:0]   _zz_mulResGroup_45_payload;
  wire       [1:0]    _zz_mulResGroup_45_payload_1;
  wire       [8:0]    _zz_mulResGroup_45_payload_2;
  wire       [8:0]    _zz_mulResGroup_45_payload_3;
  wire       [8:0]    _zz_mulResGroup_45_payload_4;
  wire       [12:0]   _zz_mulResGroup_46_payload;
  wire       [3:0]    _zz_mulResGroup_46_payload_1;
  wire       [8:0]    _zz_mulResGroup_46_payload_2;
  wire       [8:0]    _zz_mulResGroup_46_payload_3;
  wire       [8:0]    _zz_mulResGroup_46_payload_4;
  wire       [13:0]   _zz_mulResGroup_47_payload;
  wire       [4:0]    _zz_mulResGroup_47_payload_1;
  wire       [8:0]    _zz_mulResGroup_47_payload_2;
  wire       [8:0]    _zz_mulResGroup_47_payload_3;
  wire       [8:0]    _zz_mulResGroup_47_payload_4;
  wire       [13:0]   _zz_mulResGroup_48_payload;
  wire       [4:0]    _zz_mulResGroup_48_payload_1;
  wire       [8:0]    _zz_mulResGroup_48_payload_2;
  wire       [8:0]    _zz_mulResGroup_48_payload_3;
  wire       [8:0]    _zz_mulResGroup_48_payload_4;
  wire       [13:0]   _zz_mulResGroup_49_payload;
  wire       [4:0]    _zz_mulResGroup_49_payload_1;
  wire       [8:0]    _zz_mulResGroup_49_payload_2;
  wire       [8:0]    _zz_mulResGroup_49_payload_3;
  wire       [8:0]    _zz_mulResGroup_49_payload_4;
  wire       [12:0]   _zz_mulResGroup_50_payload;
  wire       [3:0]    _zz_mulResGroup_50_payload_1;
  wire       [8:0]    _zz_mulResGroup_50_payload_2;
  wire       [8:0]    _zz_mulResGroup_50_payload_3;
  wire       [8:0]    _zz_mulResGroup_50_payload_4;
  wire       [8:0]    _zz_mulResGroup_51_payload;
  wire       [12:0]   _zz_mulResGroup_52_payload;
  wire       [3:0]    _zz_mulResGroup_52_payload_1;
  wire       [8:0]    _zz_mulResGroup_52_payload_2;
  wire       [8:0]    _zz_mulResGroup_52_payload_3;
  wire       [8:0]    _zz_mulResGroup_52_payload_4;
  wire       [13:0]   _zz_mulResGroup_53_payload;
  wire       [4:0]    _zz_mulResGroup_53_payload_1;
  wire       [8:0]    _zz_mulResGroup_53_payload_2;
  wire       [8:0]    _zz_mulResGroup_53_payload_3;
  wire       [8:0]    _zz_mulResGroup_53_payload_4;
  wire       [13:0]   _zz_mulResGroup_54_payload;
  wire       [4:0]    _zz_mulResGroup_54_payload_1;
  wire       [8:0]    _zz_mulResGroup_54_payload_2;
  wire       [8:0]    _zz_mulResGroup_54_payload_3;
  wire       [8:0]    _zz_mulResGroup_54_payload_4;
  wire       [14:0]   _zz_mulResGroup_55_payload;
  wire       [5:0]    _zz_mulResGroup_55_payload_1;
  wire       [8:0]    _zz_mulResGroup_55_payload_2;
  wire       [8:0]    _zz_mulResGroup_55_payload_3;
  wire       [8:0]    _zz_mulResGroup_55_payload_4;
  wire       [13:0]   _zz_mulResGroup_56_payload;
  wire       [4:0]    _zz_mulResGroup_56_payload_1;
  wire       [8:0]    _zz_mulResGroup_56_payload_2;
  wire       [8:0]    _zz_mulResGroup_56_payload_3;
  wire       [8:0]    _zz_mulResGroup_56_payload_4;
  wire       [11:0]   _zz_mulResGroup_57_payload;
  wire       [2:0]    _zz_mulResGroup_57_payload_1;
  wire       [8:0]    _zz_mulResGroup_57_payload_2;
  wire       [8:0]    _zz_mulResGroup_57_payload_3;
  wire       [8:0]    _zz_mulResGroup_57_payload_4;
  wire       [13:0]   _zz_mulResGroup_58_payload;
  wire       [4:0]    _zz_mulResGroup_58_payload_1;
  wire       [8:0]    _zz_mulResGroup_58_payload_2;
  wire       [8:0]    _zz_mulResGroup_58_payload_3;
  wire       [8:0]    _zz_mulResGroup_58_payload_4;
  wire       [14:0]   _zz_mulResGroup_59_payload;
  wire       [5:0]    _zz_mulResGroup_59_payload_1;
  wire       [8:0]    _zz_mulResGroup_59_payload_2;
  wire       [8:0]    _zz_mulResGroup_59_payload_3;
  wire       [8:0]    _zz_mulResGroup_59_payload_4;
  wire       [15:0]   _zz_mulResGroup_60_payload;
  wire       [6:0]    _zz_mulResGroup_60_payload_1;
  wire       [8:0]    _zz_mulResGroup_60_payload_2;
  wire       [8:0]    _zz_mulResGroup_60_payload_3;
  wire       [8:0]    _zz_mulResGroup_60_payload_4;
  wire       [15:0]   _zz_mulResGroup_61_payload;
  wire       [6:0]    _zz_mulResGroup_61_payload_1;
  wire       [8:0]    _zz_mulResGroup_61_payload_2;
  wire       [8:0]    _zz_mulResGroup_61_payload_3;
  wire       [8:0]    _zz_mulResGroup_61_payload_4;
  wire       [16:0]   _zz_mulResGroup_62_payload;
  wire       [7:0]    _zz_mulResGroup_62_payload_1;
  wire       [8:0]    _zz_mulResGroup_62_payload_2;
  wire       [8:0]    _zz_mulResGroup_62_payload_3;
  wire       [8:0]    _zz_mulResGroup_62_payload_4;
  wire       [16:0]   _zz_mulResGroup_63_payload;
  wire       [7:0]    _zz_mulResGroup_63_payload_1;
  wire       [8:0]    _zz_mulResGroup_63_payload_2;
  wire       [8:0]    _zz_mulResGroup_63_payload_3;
  wire       [8:0]    _zz_mulResGroup_63_payload_4;
  wire                _zz_mulResVec_valid;
  wire                _zz_mulResVec_valid_1;
  wire                _zz_mulResVec_valid_2;
  wire       [21:0]   _zz_mulResVec_translated_payload;
  wire       [21:0]   _zz_mulResVec_translated_payload_1;
  wire       [21:0]   _zz_mulResVec_translated_payload_2;
  wire       [21:0]   _zz_mulResVec_translated_payload_3;
  wire       [21:0]   _zz_mulResVec_translated_payload_4;
  wire       [21:0]   _zz_mulResVec_translated_payload_5;
  wire       [21:0]   _zz_mulResVec_translated_payload_6;
  wire       [21:0]   _zz_mulResVec_translated_payload_7;
  wire       [21:0]   _zz_mulResVec_translated_payload_8;
  wire       [21:0]   _zz_mulResVec_translated_payload_9;
  wire       [21:0]   _zz_mulResVec_translated_payload_10;
  wire       [21:0]   _zz_mulResVec_translated_payload_11;
  wire       [21:0]   _zz_mulResVec_translated_payload_12;
  wire       [21:0]   _zz_mulResVec_translated_payload_13;
  wire       [21:0]   _zz_mulResVec_translated_payload_14;
  wire       [21:0]   _zz_mulResVec_translated_payload_15;
  wire       [21:0]   _zz_mulResVec_translated_payload_16;
  wire       [21:0]   _zz_mulResVec_translated_payload_17;
  wire       [21:0]   _zz_mulResVec_translated_payload_18;
  wire       [21:0]   _zz_mulResVec_translated_payload_19;
  wire       [21:0]   _zz_mulResVec_translated_payload_20;
  wire       [21:0]   _zz_mulResVec_translated_payload_21;
  wire       [21:0]   _zz_mulResVec_translated_payload_22;
  wire       [21:0]   _zz_mulResVec_translated_payload_23;
  wire       [21:0]   _zz_mulResVec_translated_payload_24;
  wire       [21:0]   _zz_mulResVec_translated_payload_25;
  wire       [21:0]   _zz_mulResVec_translated_payload_26;
  wire       [21:0]   _zz_mulResVec_translated_payload_27;
  wire       [21:0]   _zz_mulResVec_translated_payload_28;
  wire       [21:0]   _zz_mulResVec_translated_payload_29;
  wire       [21:0]   _zz_mulResVec_translated_payload_30;
  wire       [21:0]   _zz_mulResVec_translated_payload_31;
  wire       [21:0]   _zz_mulResVec_translated_payload_32;
  wire       [21:0]   _zz_mulResVec_translated_payload_33;
  wire       [21:0]   _zz_mulResVec_translated_payload_34;
  wire       [21:0]   _zz_mulResVec_translated_payload_35;
  wire       [21:0]   _zz_mulResVec_translated_payload_36;
  wire       [21:0]   _zz_mulResVec_translated_payload_37;
  wire       [21:0]   _zz_mulResVec_translated_payload_38;
  wire       [21:0]   _zz_mulResVec_translated_payload_39;
  wire       [21:0]   _zz_mulResVec_translated_payload_40;
  wire       [21:0]   _zz_mulResVec_translated_payload_41;
  wire       [21:0]   _zz_mulResVec_translated_payload_42;
  wire       [21:0]   _zz_mulResVec_translated_payload_43;
  wire       [21:0]   _zz_mulResVec_translated_payload_44;
  wire       [21:0]   _zz_mulResVec_translated_payload_45;
  wire       [21:0]   _zz_mulResVec_translated_payload_46;
  wire       [21:0]   _zz_mulResVec_translated_payload_47;
  wire       [21:0]   _zz_mulResVec_translated_payload_48;
  wire       [21:0]   _zz_mulResVec_translated_payload_49;
  wire       [21:0]   _zz_mulResVec_translated_payload_50;
  wire       [21:0]   _zz_mulResVec_translated_payload_51;
  wire       [21:0]   _zz_mulResVec_translated_payload_52;
  wire       [21:0]   _zz_mulResVec_translated_payload_53;
  wire       [21:0]   _zz_mulResVec_translated_payload_54;
  wire       [21:0]   _zz_mulResVec_translated_payload_55;
  wire       [21:0]   _zz_mulResVec_translated_payload_56;
  wire       [21:0]   _zz_mulResVec_translated_payload_57;
  wire       [21:0]   _zz_mulResVec_translated_payload_58;
  wire       [21:0]   _zz_mulResVec_translated_payload_59;
  wire       [21:0]   _zz_mulResVec_translated_payload_60;
  wire       [21:0]   _zz_mulResVec_translated_payload_61;
  wire                inputAll_0_valid;
  wire                inputAll_0_ready;
  wire       [7:0]    inputAll_0_payload;
  wire                inputAll_1_valid;
  wire                inputAll_1_ready;
  wire       [7:0]    inputAll_1_payload;
  wire                inputAll_2_valid;
  wire                inputAll_2_ready;
  wire       [7:0]    inputAll_2_payload;
  wire                inputAll_3_valid;
  wire                inputAll_3_ready;
  wire       [7:0]    inputAll_3_payload;
  wire                inputAll_4_valid;
  wire                inputAll_4_ready;
  wire       [7:0]    inputAll_4_payload;
  wire                inputAll_5_valid;
  wire                inputAll_5_ready;
  wire       [7:0]    inputAll_5_payload;
  wire                inputAll_6_valid;
  wire                inputAll_6_ready;
  wire       [7:0]    inputAll_6_payload;
  wire                inputAll_7_valid;
  wire                inputAll_7_ready;
  wire       [7:0]    inputAll_7_payload;
  wire                inputAll_8_valid;
  wire                inputAll_8_ready;
  wire       [7:0]    inputAll_8_payload;
  wire                inputAll_9_valid;
  wire                inputAll_9_ready;
  wire       [7:0]    inputAll_9_payload;
  wire                inputAll_10_valid;
  wire                inputAll_10_ready;
  wire       [7:0]    inputAll_10_payload;
  wire                inputAll_11_valid;
  wire                inputAll_11_ready;
  wire       [7:0]    inputAll_11_payload;
  wire                inputAll_12_valid;
  wire                inputAll_12_ready;
  wire       [7:0]    inputAll_12_payload;
  wire                inputAll_13_valid;
  wire                inputAll_13_ready;
  wire       [7:0]    inputAll_13_payload;
  wire                inputAll_14_valid;
  wire                inputAll_14_ready;
  wire       [7:0]    inputAll_14_payload;
  wire                inputAll_15_valid;
  wire                inputAll_15_ready;
  wire       [7:0]    inputAll_15_payload;
  wire                inputAll_16_valid;
  wire                inputAll_16_ready;
  wire       [7:0]    inputAll_16_payload;
  wire                inputAll_17_valid;
  wire                inputAll_17_ready;
  wire       [7:0]    inputAll_17_payload;
  wire                inputAll_18_valid;
  wire                inputAll_18_ready;
  wire       [7:0]    inputAll_18_payload;
  wire                inputAll_19_valid;
  wire                inputAll_19_ready;
  wire       [7:0]    inputAll_19_payload;
  wire                inputAll_20_valid;
  wire                inputAll_20_ready;
  wire       [7:0]    inputAll_20_payload;
  wire                inputAll_21_valid;
  wire                inputAll_21_ready;
  wire       [7:0]    inputAll_21_payload;
  wire                inputAll_22_valid;
  wire                inputAll_22_ready;
  wire       [7:0]    inputAll_22_payload;
  wire                inputAll_23_valid;
  wire                inputAll_23_ready;
  wire       [7:0]    inputAll_23_payload;
  wire                inputAll_24_valid;
  wire                inputAll_24_ready;
  wire       [7:0]    inputAll_24_payload;
  wire                inputAll_25_valid;
  wire                inputAll_25_ready;
  wire       [7:0]    inputAll_25_payload;
  wire                inputAll_26_valid;
  wire                inputAll_26_ready;
  wire       [7:0]    inputAll_26_payload;
  wire                inputAll_27_valid;
  wire                inputAll_27_ready;
  wire       [7:0]    inputAll_27_payload;
  wire                inputAll_28_valid;
  wire                inputAll_28_ready;
  wire       [7:0]    inputAll_28_payload;
  wire                inputAll_29_valid;
  wire                inputAll_29_ready;
  wire       [7:0]    inputAll_29_payload;
  wire                inputAll_30_valid;
  wire                inputAll_30_ready;
  wire       [7:0]    inputAll_30_payload;
  wire                inputAll_31_valid;
  wire                inputAll_31_ready;
  wire       [7:0]    inputAll_31_payload;
  wire                inputAll_32_valid;
  wire                inputAll_32_ready;
  wire       [7:0]    inputAll_32_payload;
  wire                inputAll_33_valid;
  wire                inputAll_33_ready;
  wire       [7:0]    inputAll_33_payload;
  wire                inputAll_34_valid;
  wire                inputAll_34_ready;
  wire       [7:0]    inputAll_34_payload;
  wire                inputAll_35_valid;
  wire                inputAll_35_ready;
  wire       [7:0]    inputAll_35_payload;
  wire                inputAll_36_valid;
  wire                inputAll_36_ready;
  wire       [7:0]    inputAll_36_payload;
  wire                inputAll_37_valid;
  wire                inputAll_37_ready;
  wire       [7:0]    inputAll_37_payload;
  wire                inputAll_38_valid;
  wire                inputAll_38_ready;
  wire       [7:0]    inputAll_38_payload;
  wire                inputAll_39_valid;
  wire                inputAll_39_ready;
  wire       [7:0]    inputAll_39_payload;
  wire                inputAll_40_valid;
  wire                inputAll_40_ready;
  wire       [7:0]    inputAll_40_payload;
  wire                inputAll_41_valid;
  wire                inputAll_41_ready;
  wire       [7:0]    inputAll_41_payload;
  wire                inputAll_42_valid;
  wire                inputAll_42_ready;
  wire       [7:0]    inputAll_42_payload;
  wire                inputAll_43_valid;
  wire                inputAll_43_ready;
  wire       [7:0]    inputAll_43_payload;
  wire                inputAll_44_valid;
  wire                inputAll_44_ready;
  wire       [7:0]    inputAll_44_payload;
  wire                inputAll_45_valid;
  wire                inputAll_45_ready;
  wire       [7:0]    inputAll_45_payload;
  wire                inputAll_46_valid;
  wire                inputAll_46_ready;
  wire       [7:0]    inputAll_46_payload;
  wire                inputAll_47_valid;
  wire                inputAll_47_ready;
  wire       [7:0]    inputAll_47_payload;
  wire                inputAll_48_valid;
  wire                inputAll_48_ready;
  wire       [7:0]    inputAll_48_payload;
  wire                inputAll_49_valid;
  wire                inputAll_49_ready;
  wire       [7:0]    inputAll_49_payload;
  wire                inputAll_50_valid;
  wire                inputAll_50_ready;
  wire       [7:0]    inputAll_50_payload;
  wire                inputAll_51_valid;
  wire                inputAll_51_ready;
  wire       [7:0]    inputAll_51_payload;
  wire                inputAll_52_valid;
  wire                inputAll_52_ready;
  wire       [7:0]    inputAll_52_payload;
  wire                inputAll_53_valid;
  wire                inputAll_53_ready;
  wire       [7:0]    inputAll_53_payload;
  wire                inputAll_54_valid;
  wire                inputAll_54_ready;
  wire       [7:0]    inputAll_54_payload;
  wire                inputAll_55_valid;
  wire                inputAll_55_ready;
  wire       [7:0]    inputAll_55_payload;
  wire                inputAll_56_valid;
  wire                inputAll_56_ready;
  wire       [7:0]    inputAll_56_payload;
  wire                inputAll_57_valid;
  wire                inputAll_57_ready;
  wire       [7:0]    inputAll_57_payload;
  wire                inputAll_58_valid;
  wire                inputAll_58_ready;
  wire       [7:0]    inputAll_58_payload;
  wire                inputAll_59_valid;
  wire                inputAll_59_ready;
  wire       [7:0]    inputAll_59_payload;
  wire                inputAll_60_valid;
  wire                inputAll_60_ready;
  wire       [7:0]    inputAll_60_payload;
  wire                inputAll_61_valid;
  wire                inputAll_61_ready;
  wire       [7:0]    inputAll_61_payload;
  wire                inputAll_62_valid;
  wire                inputAll_62_ready;
  wire       [7:0]    inputAll_62_payload;
  wire                inputAll_63_valid;
  wire                inputAll_63_ready;
  wire       [7:0]    inputAll_63_payload;
  wire                inputAll_64_valid;
  wire                inputAll_64_ready;
  wire       [7:0]    inputAll_64_payload;
  wire                inputAll_65_valid;
  wire                inputAll_65_ready;
  wire       [7:0]    inputAll_65_payload;
  wire                inputAll_66_valid;
  wire                inputAll_66_ready;
  wire       [7:0]    inputAll_66_payload;
  wire                inputAll_67_valid;
  wire                inputAll_67_ready;
  wire       [7:0]    inputAll_67_payload;
  wire                inputAll_68_valid;
  wire                inputAll_68_ready;
  wire       [7:0]    inputAll_68_payload;
  wire                inputAll_69_valid;
  wire                inputAll_69_ready;
  wire       [7:0]    inputAll_69_payload;
  wire                inputAll_70_valid;
  wire                inputAll_70_ready;
  wire       [7:0]    inputAll_70_payload;
  wire                inputAll_71_valid;
  wire                inputAll_71_ready;
  wire       [7:0]    inputAll_71_payload;
  wire                inputAll_72_valid;
  wire                inputAll_72_ready;
  wire       [7:0]    inputAll_72_payload;
  wire                inputAll_73_valid;
  wire                inputAll_73_ready;
  wire       [7:0]    inputAll_73_payload;
  wire                inputAll_74_valid;
  wire                inputAll_74_ready;
  wire       [7:0]    inputAll_74_payload;
  wire                inputAll_75_valid;
  wire                inputAll_75_ready;
  wire       [7:0]    inputAll_75_payload;
  wire                inputAll_76_valid;
  wire                inputAll_76_ready;
  wire       [7:0]    inputAll_76_payload;
  wire                inputAll_77_valid;
  wire                inputAll_77_ready;
  wire       [7:0]    inputAll_77_payload;
  wire                inputAll_78_valid;
  wire                inputAll_78_ready;
  wire       [7:0]    inputAll_78_payload;
  wire                inputAll_79_valid;
  wire                inputAll_79_ready;
  wire       [7:0]    inputAll_79_payload;
  wire                inputAll_80_valid;
  wire                inputAll_80_ready;
  wire       [7:0]    inputAll_80_payload;
  wire                inputAll_81_valid;
  wire                inputAll_81_ready;
  wire       [7:0]    inputAll_81_payload;
  wire                inputAll_82_valid;
  wire                inputAll_82_ready;
  wire       [7:0]    inputAll_82_payload;
  wire                inputAll_83_valid;
  wire                inputAll_83_ready;
  wire       [7:0]    inputAll_83_payload;
  wire                inputAll_84_valid;
  wire                inputAll_84_ready;
  wire       [7:0]    inputAll_84_payload;
  wire                inputAll_85_valid;
  wire                inputAll_85_ready;
  wire       [7:0]    inputAll_85_payload;
  wire                inputAll_86_valid;
  wire                inputAll_86_ready;
  wire       [7:0]    inputAll_86_payload;
  wire                inputAll_87_valid;
  wire                inputAll_87_ready;
  wire       [7:0]    inputAll_87_payload;
  wire                inputAll_88_valid;
  wire                inputAll_88_ready;
  wire       [7:0]    inputAll_88_payload;
  wire                inputAll_89_valid;
  wire                inputAll_89_ready;
  wire       [7:0]    inputAll_89_payload;
  wire                inputAll_90_valid;
  wire                inputAll_90_ready;
  wire       [7:0]    inputAll_90_payload;
  wire                inputAll_91_valid;
  wire                inputAll_91_ready;
  wire       [7:0]    inputAll_91_payload;
  wire                inputAll_92_valid;
  wire                inputAll_92_ready;
  wire       [7:0]    inputAll_92_payload;
  wire                inputAll_93_valid;
  wire                inputAll_93_ready;
  wire       [7:0]    inputAll_93_payload;
  wire                inputAll_94_valid;
  wire                inputAll_94_ready;
  wire       [7:0]    inputAll_94_payload;
  wire                inputAll_95_valid;
  wire                inputAll_95_ready;
  wire       [7:0]    inputAll_95_payload;
  wire                inputAll_96_valid;
  wire                inputAll_96_ready;
  wire       [7:0]    inputAll_96_payload;
  wire                inputAll_97_valid;
  wire                inputAll_97_ready;
  wire       [7:0]    inputAll_97_payload;
  wire                inputAll_98_valid;
  wire                inputAll_98_ready;
  wire       [7:0]    inputAll_98_payload;
  wire                inputAll_99_valid;
  wire                inputAll_99_ready;
  wire       [7:0]    inputAll_99_payload;
  wire                inputAll_100_valid;
  wire                inputAll_100_ready;
  wire       [7:0]    inputAll_100_payload;
  wire                inputAll_101_valid;
  wire                inputAll_101_ready;
  wire       [7:0]    inputAll_101_payload;
  wire                inputAll_102_valid;
  wire                inputAll_102_ready;
  wire       [7:0]    inputAll_102_payload;
  wire                inputAll_103_valid;
  wire                inputAll_103_ready;
  wire       [7:0]    inputAll_103_payload;
  wire                inputAll_104_valid;
  wire                inputAll_104_ready;
  wire       [7:0]    inputAll_104_payload;
  wire                inputAll_105_valid;
  wire                inputAll_105_ready;
  wire       [7:0]    inputAll_105_payload;
  wire                inputAll_106_valid;
  wire                inputAll_106_ready;
  wire       [7:0]    inputAll_106_payload;
  wire                inputAll_107_valid;
  wire                inputAll_107_ready;
  wire       [7:0]    inputAll_107_payload;
  wire                inputAll_108_valid;
  wire                inputAll_108_ready;
  wire       [7:0]    inputAll_108_payload;
  wire                inputAll_109_valid;
  wire                inputAll_109_ready;
  wire       [7:0]    inputAll_109_payload;
  wire                inputAll_110_valid;
  wire                inputAll_110_ready;
  wire       [7:0]    inputAll_110_payload;
  wire                inputAll_111_valid;
  wire                inputAll_111_ready;
  wire       [7:0]    inputAll_111_payload;
  wire                inputAll_112_valid;
  wire                inputAll_112_ready;
  wire       [7:0]    inputAll_112_payload;
  wire                inputAll_113_valid;
  wire                inputAll_113_ready;
  wire       [7:0]    inputAll_113_payload;
  wire                inputAll_114_valid;
  wire                inputAll_114_ready;
  wire       [7:0]    inputAll_114_payload;
  wire                inputAll_115_valid;
  wire                inputAll_115_ready;
  wire       [7:0]    inputAll_115_payload;
  wire                inputAll_116_valid;
  wire                inputAll_116_ready;
  wire       [7:0]    inputAll_116_payload;
  wire                inputAll_117_valid;
  wire                inputAll_117_ready;
  wire       [7:0]    inputAll_117_payload;
  wire                inputAll_118_valid;
  wire                inputAll_118_ready;
  wire       [7:0]    inputAll_118_payload;
  wire                inputAll_119_valid;
  wire                inputAll_119_ready;
  wire       [7:0]    inputAll_119_payload;
  wire                inputAll_120_valid;
  wire                inputAll_120_ready;
  wire       [7:0]    inputAll_120_payload;
  wire                inputAll_121_valid;
  wire                inputAll_121_ready;
  wire       [7:0]    inputAll_121_payload;
  wire                inputAll_122_valid;
  wire                inputAll_122_ready;
  wire       [7:0]    inputAll_122_payload;
  wire                inputAll_123_valid;
  wire                inputAll_123_ready;
  wire       [7:0]    inputAll_123_payload;
  wire                inputAll_124_valid;
  wire                inputAll_124_ready;
  wire       [7:0]    inputAll_124_payload;
  wire                inputAll_125_valid;
  wire                inputAll_125_ready;
  wire       [7:0]    inputAll_125_payload;
  wire                inputAll_126_valid;
  wire                inputAll_126_ready;
  wire       [7:0]    inputAll_126_payload;
  wire                inputAll_127_valid;
  wire                inputAll_127_ready;
  wire       [7:0]    inputAll_127_payload;
  wire                inputAll_0_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_0_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_0_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_0_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_0_fork_io_outputs_1_rData;
  wire                when_Stream_l342;
  wire                inputAll_1_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_1_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_1_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_1_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_1_fork_io_outputs_1_rData;
  wire                when_Stream_l342_1;
  wire                inputAll_2_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_2_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_2_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_2_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_2_fork_io_outputs_1_rData;
  wire                when_Stream_l342_2;
  wire                inputAll_3_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_3_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_3_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_3_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_3_fork_io_outputs_1_rData;
  wire                when_Stream_l342_3;
  wire                inputAll_4_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_4_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_4_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_4_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_4_fork_io_outputs_1_rData;
  wire                when_Stream_l342_4;
  wire                inputAll_5_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_5_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_5_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_5_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_5_fork_io_outputs_1_rData;
  wire                when_Stream_l342_5;
  wire                inputAll_6_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_6_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_6_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_6_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_6_fork_io_outputs_1_rData;
  wire                when_Stream_l342_6;
  wire                inputAll_7_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_7_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_7_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_7_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_7_fork_io_outputs_1_rData;
  wire                when_Stream_l342_7;
  wire                inputAll_8_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_8_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_8_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_8_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_8_fork_io_outputs_1_rData;
  wire                when_Stream_l342_8;
  wire                inputAll_9_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_9_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_9_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_9_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_9_fork_io_outputs_1_rData;
  wire                when_Stream_l342_9;
  wire                inputAll_10_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_10_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_10_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_10_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_10_fork_io_outputs_1_rData;
  wire                when_Stream_l342_10;
  wire                inputAll_11_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_11_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_11_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_11_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_11_fork_io_outputs_1_rData;
  wire                when_Stream_l342_11;
  wire                inputAll_12_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_12_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_12_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_12_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_12_fork_io_outputs_1_rData;
  wire                when_Stream_l342_12;
  wire                inputAll_13_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_13_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_13_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_13_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_13_fork_io_outputs_1_rData;
  wire                when_Stream_l342_13;
  wire                inputAll_14_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_14_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_14_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_14_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_14_fork_io_outputs_1_rData;
  wire                when_Stream_l342_14;
  wire                inputAll_15_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_15_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_15_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_15_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_15_fork_io_outputs_1_rData;
  wire                when_Stream_l342_15;
  wire                inputAll_16_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_16_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_16_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_16_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_16_fork_io_outputs_1_rData;
  wire                when_Stream_l342_16;
  wire                inputAll_17_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_17_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_17_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_17_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_17_fork_io_outputs_1_rData;
  wire                when_Stream_l342_17;
  wire                inputAll_18_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_18_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_18_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_18_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_18_fork_io_outputs_1_rData;
  wire                when_Stream_l342_18;
  wire                inputAll_19_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_19_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_19_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_19_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_19_fork_io_outputs_1_rData;
  wire                when_Stream_l342_19;
  wire                inputAll_20_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_20_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_20_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_20_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_20_fork_io_outputs_1_rData;
  wire                when_Stream_l342_20;
  wire                inputAll_21_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_21_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_21_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_21_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_21_fork_io_outputs_1_rData;
  wire                when_Stream_l342_21;
  wire                inputAll_22_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_22_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_22_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_22_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_22_fork_io_outputs_1_rData;
  wire                when_Stream_l342_22;
  wire                inputAll_23_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_23_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_23_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_23_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_23_fork_io_outputs_1_rData;
  wire                when_Stream_l342_23;
  wire                inputAll_24_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_24_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_24_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_24_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_24_fork_io_outputs_1_rData;
  wire                when_Stream_l342_24;
  wire                inputAll_25_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_25_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_25_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_25_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_25_fork_io_outputs_1_rData;
  wire                when_Stream_l342_25;
  wire                inputAll_26_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_26_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_26_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_26_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_26_fork_io_outputs_1_rData;
  wire                when_Stream_l342_26;
  wire                inputAll_27_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_27_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_27_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_27_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_27_fork_io_outputs_1_rData;
  wire                when_Stream_l342_27;
  wire                inputAll_28_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_28_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_28_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_28_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_28_fork_io_outputs_1_rData;
  wire                when_Stream_l342_28;
  wire                inputAll_29_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_29_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_29_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_29_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_29_fork_io_outputs_1_rData;
  wire                when_Stream_l342_29;
  wire                inputAll_30_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_30_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_30_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_30_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_30_fork_io_outputs_1_rData;
  wire                when_Stream_l342_30;
  wire                inputAll_31_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_31_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_31_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_31_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_31_fork_io_outputs_1_rData;
  wire                when_Stream_l342_31;
  wire                inputAll_32_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_32_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_32_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_32_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_32_fork_io_outputs_1_rData;
  wire                when_Stream_l342_32;
  wire                inputAll_33_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_33_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_33_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_33_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_33_fork_io_outputs_1_rData;
  wire                when_Stream_l342_33;
  wire                inputAll_34_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_34_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_34_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_34_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_34_fork_io_outputs_1_rData;
  wire                when_Stream_l342_34;
  wire                inputAll_35_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_35_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_35_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_35_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_35_fork_io_outputs_1_rData;
  wire                when_Stream_l342_35;
  wire                inputAll_36_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_36_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_36_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_36_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_36_fork_io_outputs_1_rData;
  wire                when_Stream_l342_36;
  wire                inputAll_37_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_37_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_37_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_37_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_37_fork_io_outputs_1_rData;
  wire                when_Stream_l342_37;
  wire                inputAll_38_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_38_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_38_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_38_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_38_fork_io_outputs_1_rData;
  wire                when_Stream_l342_38;
  wire                inputAll_39_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_39_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_39_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_39_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_39_fork_io_outputs_1_rData;
  wire                when_Stream_l342_39;
  wire                inputAll_40_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_40_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_40_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_40_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_40_fork_io_outputs_1_rData;
  wire                when_Stream_l342_40;
  wire                inputAll_41_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_41_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_41_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_41_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_41_fork_io_outputs_1_rData;
  wire                when_Stream_l342_41;
  wire                inputAll_42_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_42_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_42_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_42_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_42_fork_io_outputs_1_rData;
  wire                when_Stream_l342_42;
  wire                inputAll_43_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_43_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_43_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_43_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_43_fork_io_outputs_1_rData;
  wire                when_Stream_l342_43;
  wire                inputAll_44_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_44_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_44_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_44_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_44_fork_io_outputs_1_rData;
  wire                when_Stream_l342_44;
  wire                inputAll_45_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_45_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_45_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_45_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_45_fork_io_outputs_1_rData;
  wire                when_Stream_l342_45;
  wire                inputAll_46_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_46_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_46_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_46_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_46_fork_io_outputs_1_rData;
  wire                when_Stream_l342_46;
  wire                inputAll_47_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_47_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_47_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_47_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_47_fork_io_outputs_1_rData;
  wire                when_Stream_l342_47;
  wire                inputAll_48_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_48_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_48_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_48_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_48_fork_io_outputs_1_rData;
  wire                when_Stream_l342_48;
  wire                inputAll_49_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_49_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_49_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_49_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_49_fork_io_outputs_1_rData;
  wire                when_Stream_l342_49;
  wire                inputAll_50_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_50_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_50_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_50_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_50_fork_io_outputs_1_rData;
  wire                when_Stream_l342_50;
  wire                inputAll_51_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_51_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_51_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_51_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_51_fork_io_outputs_1_rData;
  wire                when_Stream_l342_51;
  wire                inputAll_52_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_52_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_52_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_52_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_52_fork_io_outputs_1_rData;
  wire                when_Stream_l342_52;
  wire                inputAll_53_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_53_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_53_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_53_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_53_fork_io_outputs_1_rData;
  wire                when_Stream_l342_53;
  wire                inputAll_54_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_54_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_54_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_54_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_54_fork_io_outputs_1_rData;
  wire                when_Stream_l342_54;
  wire                inputAll_55_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_55_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_55_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_55_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_55_fork_io_outputs_1_rData;
  wire                when_Stream_l342_55;
  wire                inputAll_56_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_56_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_56_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_56_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_56_fork_io_outputs_1_rData;
  wire                when_Stream_l342_56;
  wire                inputAll_57_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_57_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_57_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_57_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_57_fork_io_outputs_1_rData;
  wire                when_Stream_l342_57;
  wire                inputAll_58_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_58_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_58_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_58_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_58_fork_io_outputs_1_rData;
  wire                when_Stream_l342_58;
  wire                inputAll_59_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_59_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_59_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_59_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_59_fork_io_outputs_1_rData;
  wire                when_Stream_l342_59;
  wire                inputAll_60_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_60_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_60_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_60_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_60_fork_io_outputs_1_rData;
  wire                when_Stream_l342_60;
  wire                inputAll_61_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_61_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_61_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_61_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_61_fork_io_outputs_1_rData;
  wire                when_Stream_l342_61;
  wire                inputAll_62_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_62_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_62_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_62_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_62_fork_io_outputs_1_rData;
  wire                when_Stream_l342_62;
  wire                inputAll_63_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_63_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_63_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_63_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_63_fork_io_outputs_1_rData;
  wire                when_Stream_l342_63;
  wire                inputAll_64_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_64_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_64_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_64_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_64_fork_io_outputs_1_rData;
  wire                when_Stream_l342_64;
  wire                inputAll_65_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_65_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_65_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_65_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_65_fork_io_outputs_1_rData;
  wire                when_Stream_l342_65;
  wire                inputAll_66_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_66_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_66_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_66_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_66_fork_io_outputs_1_rData;
  wire                when_Stream_l342_66;
  wire                inputAll_67_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_67_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_67_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_67_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_67_fork_io_outputs_1_rData;
  wire                when_Stream_l342_67;
  wire                inputAll_68_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_68_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_68_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_68_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_68_fork_io_outputs_1_rData;
  wire                when_Stream_l342_68;
  wire                inputAll_69_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_69_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_69_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_69_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_69_fork_io_outputs_1_rData;
  wire                when_Stream_l342_69;
  wire                inputAll_70_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_70_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_70_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_70_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_70_fork_io_outputs_1_rData;
  wire                when_Stream_l342_70;
  wire                inputAll_71_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_71_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_71_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_71_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_71_fork_io_outputs_1_rData;
  wire                when_Stream_l342_71;
  wire                inputAll_72_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_72_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_72_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_72_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_72_fork_io_outputs_1_rData;
  wire                when_Stream_l342_72;
  wire                inputAll_73_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_73_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_73_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_73_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_73_fork_io_outputs_1_rData;
  wire                when_Stream_l342_73;
  wire                inputAll_74_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_74_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_74_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_74_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_74_fork_io_outputs_1_rData;
  wire                when_Stream_l342_74;
  wire                inputAll_75_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_75_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_75_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_75_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_75_fork_io_outputs_1_rData;
  wire                when_Stream_l342_75;
  wire                inputAll_76_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_76_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_76_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_76_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_76_fork_io_outputs_1_rData;
  wire                when_Stream_l342_76;
  wire                inputAll_77_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_77_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_77_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_77_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_77_fork_io_outputs_1_rData;
  wire                when_Stream_l342_77;
  wire                inputAll_78_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_78_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_78_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_78_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_78_fork_io_outputs_1_rData;
  wire                when_Stream_l342_78;
  wire                inputAll_79_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_79_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_79_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_79_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_79_fork_io_outputs_1_rData;
  wire                when_Stream_l342_79;
  wire                inputAll_80_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_80_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_80_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_80_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_80_fork_io_outputs_1_rData;
  wire                when_Stream_l342_80;
  wire                inputAll_81_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_81_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_81_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_81_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_81_fork_io_outputs_1_rData;
  wire                when_Stream_l342_81;
  wire                inputAll_82_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_82_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_82_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_82_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_82_fork_io_outputs_1_rData;
  wire                when_Stream_l342_82;
  wire                inputAll_83_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_83_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_83_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_83_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_83_fork_io_outputs_1_rData;
  wire                when_Stream_l342_83;
  wire                inputAll_84_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_84_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_84_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_84_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_84_fork_io_outputs_1_rData;
  wire                when_Stream_l342_84;
  wire                inputAll_85_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_85_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_85_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_85_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_85_fork_io_outputs_1_rData;
  wire                when_Stream_l342_85;
  wire                inputAll_86_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_86_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_86_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_86_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_86_fork_io_outputs_1_rData;
  wire                when_Stream_l342_86;
  wire                inputAll_87_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_87_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_87_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_87_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_87_fork_io_outputs_1_rData;
  wire                when_Stream_l342_87;
  wire                inputAll_88_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_88_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_88_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_88_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_88_fork_io_outputs_1_rData;
  wire                when_Stream_l342_88;
  wire                inputAll_89_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_89_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_89_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_89_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_89_fork_io_outputs_1_rData;
  wire                when_Stream_l342_89;
  wire                inputAll_90_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_90_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_90_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_90_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_90_fork_io_outputs_1_rData;
  wire                when_Stream_l342_90;
  wire                inputAll_91_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_91_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_91_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_91_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_91_fork_io_outputs_1_rData;
  wire                when_Stream_l342_91;
  wire                inputAll_92_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_92_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_92_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_92_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_92_fork_io_outputs_1_rData;
  wire                when_Stream_l342_92;
  wire                inputAll_93_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_93_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_93_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_93_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_93_fork_io_outputs_1_rData;
  wire                when_Stream_l342_93;
  wire                inputAll_94_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_94_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_94_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_94_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_94_fork_io_outputs_1_rData;
  wire                when_Stream_l342_94;
  wire                inputAll_95_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_95_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_95_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_95_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_95_fork_io_outputs_1_rData;
  wire                when_Stream_l342_95;
  wire                inputAll_96_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_96_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_96_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_96_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_96_fork_io_outputs_1_rData;
  wire                when_Stream_l342_96;
  wire                inputAll_97_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_97_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_97_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_97_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_97_fork_io_outputs_1_rData;
  wire                when_Stream_l342_97;
  wire                inputAll_98_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_98_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_98_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_98_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_98_fork_io_outputs_1_rData;
  wire                when_Stream_l342_98;
  wire                inputAll_99_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_99_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_99_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_99_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_99_fork_io_outputs_1_rData;
  wire                when_Stream_l342_99;
  wire                inputAll_100_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_100_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_100_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_100_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_100_fork_io_outputs_1_rData;
  wire                when_Stream_l342_100;
  wire                inputAll_101_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_101_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_101_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_101_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_101_fork_io_outputs_1_rData;
  wire                when_Stream_l342_101;
  wire                inputAll_102_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_102_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_102_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_102_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_102_fork_io_outputs_1_rData;
  wire                when_Stream_l342_102;
  wire                inputAll_103_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_103_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_103_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_103_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_103_fork_io_outputs_1_rData;
  wire                when_Stream_l342_103;
  wire                inputAll_104_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_104_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_104_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_104_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_104_fork_io_outputs_1_rData;
  wire                when_Stream_l342_104;
  wire                inputAll_105_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_105_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_105_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_105_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_105_fork_io_outputs_1_rData;
  wire                when_Stream_l342_105;
  wire                inputAll_106_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_106_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_106_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_106_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_106_fork_io_outputs_1_rData;
  wire                when_Stream_l342_106;
  wire                inputAll_107_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_107_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_107_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_107_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_107_fork_io_outputs_1_rData;
  wire                when_Stream_l342_107;
  wire                inputAll_108_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_108_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_108_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_108_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_108_fork_io_outputs_1_rData;
  wire                when_Stream_l342_108;
  wire                inputAll_109_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_109_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_109_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_109_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_109_fork_io_outputs_1_rData;
  wire                when_Stream_l342_109;
  wire                inputAll_110_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_110_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_110_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_110_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_110_fork_io_outputs_1_rData;
  wire                when_Stream_l342_110;
  wire                inputAll_111_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_111_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_111_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_111_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_111_fork_io_outputs_1_rData;
  wire                when_Stream_l342_111;
  wire                inputAll_112_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_112_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_112_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_112_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_112_fork_io_outputs_1_rData;
  wire                when_Stream_l342_112;
  wire                inputAll_113_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_113_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_113_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_113_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_113_fork_io_outputs_1_rData;
  wire                when_Stream_l342_113;
  wire                inputAll_114_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_114_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_114_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_114_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_114_fork_io_outputs_1_rData;
  wire                when_Stream_l342_114;
  wire                inputAll_115_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_115_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_115_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_115_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_115_fork_io_outputs_1_rData;
  wire                when_Stream_l342_115;
  wire                inputAll_116_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_116_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_116_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_116_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_116_fork_io_outputs_1_rData;
  wire                when_Stream_l342_116;
  wire                inputAll_117_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_117_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_117_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_117_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_117_fork_io_outputs_1_rData;
  wire                when_Stream_l342_117;
  wire                inputAll_118_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_118_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_118_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_118_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_118_fork_io_outputs_1_rData;
  wire                when_Stream_l342_118;
  wire                inputAll_119_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_119_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_119_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_119_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_119_fork_io_outputs_1_rData;
  wire                when_Stream_l342_119;
  wire                inputAll_120_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_120_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_120_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_120_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_120_fork_io_outputs_1_rData;
  wire                when_Stream_l342_120;
  wire                inputAll_121_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_121_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_121_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_121_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_121_fork_io_outputs_1_rData;
  wire                when_Stream_l342_121;
  wire                inputAll_122_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_122_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_122_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_122_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_122_fork_io_outputs_1_rData;
  wire                when_Stream_l342_122;
  wire                inputAll_123_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_123_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_123_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_123_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_123_fork_io_outputs_1_rData;
  wire                when_Stream_l342_123;
  wire                inputAll_124_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_124_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_124_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_124_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_124_fork_io_outputs_1_rData;
  wire                when_Stream_l342_124;
  wire                inputAll_125_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_125_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_125_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_125_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_125_fork_io_outputs_1_rData;
  wire                when_Stream_l342_125;
  wire                inputAll_126_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_126_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_126_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_126_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_126_fork_io_outputs_1_rData;
  wire                when_Stream_l342_126;
  wire                inputAll_127_fork_io_outputs_1_m2sPipe_valid;
  wire                inputAll_127_fork_io_outputs_1_m2sPipe_ready;
  wire       [7:0]    inputAll_127_fork_io_outputs_1_m2sPipe_payload;
  reg                 inputAll_127_fork_io_outputs_1_rValid;
  reg        [7:0]    inputAll_127_fork_io_outputs_1_rData;
  wire                when_Stream_l342_127;
  wire                mulResGroup_0_valid;
  wire                mulResGroup_0_ready;
  wire       [21:0]   mulResGroup_0_payload;
  wire                mulResGroup_1_valid;
  wire                mulResGroup_1_ready;
  wire       [21:0]   mulResGroup_1_payload;
  wire                mulResGroup_2_valid;
  wire                mulResGroup_2_ready;
  wire       [21:0]   mulResGroup_2_payload;
  wire                mulResGroup_3_valid;
  wire                mulResGroup_3_ready;
  wire       [21:0]   mulResGroup_3_payload;
  wire                mulResGroup_4_valid;
  wire                mulResGroup_4_ready;
  wire       [21:0]   mulResGroup_4_payload;
  wire                mulResGroup_5_valid;
  wire                mulResGroup_5_ready;
  wire       [21:0]   mulResGroup_5_payload;
  wire                mulResGroup_6_valid;
  wire                mulResGroup_6_ready;
  wire       [21:0]   mulResGroup_6_payload;
  wire                mulResGroup_7_valid;
  wire                mulResGroup_7_ready;
  wire       [21:0]   mulResGroup_7_payload;
  wire                mulResGroup_8_valid;
  wire                mulResGroup_8_ready;
  wire       [21:0]   mulResGroup_8_payload;
  wire                mulResGroup_9_valid;
  wire                mulResGroup_9_ready;
  wire       [21:0]   mulResGroup_9_payload;
  wire                mulResGroup_10_valid;
  wire                mulResGroup_10_ready;
  wire       [21:0]   mulResGroup_10_payload;
  wire                mulResGroup_11_valid;
  wire                mulResGroup_11_ready;
  wire       [21:0]   mulResGroup_11_payload;
  wire                mulResGroup_12_valid;
  wire                mulResGroup_12_ready;
  wire       [21:0]   mulResGroup_12_payload;
  wire                mulResGroup_13_valid;
  wire                mulResGroup_13_ready;
  wire       [21:0]   mulResGroup_13_payload;
  wire                mulResGroup_14_valid;
  wire                mulResGroup_14_ready;
  wire       [21:0]   mulResGroup_14_payload;
  wire                mulResGroup_15_valid;
  wire                mulResGroup_15_ready;
  wire       [21:0]   mulResGroup_15_payload;
  wire                mulResGroup_16_valid;
  wire                mulResGroup_16_ready;
  wire       [21:0]   mulResGroup_16_payload;
  wire                mulResGroup_17_valid;
  wire                mulResGroup_17_ready;
  wire       [21:0]   mulResGroup_17_payload;
  wire                mulResGroup_18_valid;
  wire                mulResGroup_18_ready;
  wire       [21:0]   mulResGroup_18_payload;
  wire                mulResGroup_19_valid;
  wire                mulResGroup_19_ready;
  wire       [21:0]   mulResGroup_19_payload;
  wire                mulResGroup_20_valid;
  wire                mulResGroup_20_ready;
  wire       [21:0]   mulResGroup_20_payload;
  wire                mulResGroup_21_valid;
  wire                mulResGroup_21_ready;
  wire       [21:0]   mulResGroup_21_payload;
  wire                mulResGroup_22_valid;
  wire                mulResGroup_22_ready;
  wire       [21:0]   mulResGroup_22_payload;
  wire                mulResGroup_23_valid;
  wire                mulResGroup_23_ready;
  wire       [21:0]   mulResGroup_23_payload;
  wire                mulResGroup_24_valid;
  wire                mulResGroup_24_ready;
  wire       [21:0]   mulResGroup_24_payload;
  wire                mulResGroup_25_valid;
  wire                mulResGroup_25_ready;
  wire       [21:0]   mulResGroup_25_payload;
  wire                mulResGroup_26_valid;
  wire                mulResGroup_26_ready;
  wire       [21:0]   mulResGroup_26_payload;
  wire                mulResGroup_27_valid;
  wire                mulResGroup_27_ready;
  wire       [21:0]   mulResGroup_27_payload;
  wire                mulResGroup_28_valid;
  wire                mulResGroup_28_ready;
  wire       [21:0]   mulResGroup_28_payload;
  wire                mulResGroup_29_valid;
  wire                mulResGroup_29_ready;
  wire       [21:0]   mulResGroup_29_payload;
  wire                mulResGroup_30_valid;
  wire                mulResGroup_30_ready;
  wire       [21:0]   mulResGroup_30_payload;
  wire                mulResGroup_31_valid;
  wire                mulResGroup_31_ready;
  wire       [21:0]   mulResGroup_31_payload;
  wire                mulResGroup_32_valid;
  wire                mulResGroup_32_ready;
  wire       [21:0]   mulResGroup_32_payload;
  wire                mulResGroup_33_valid;
  wire                mulResGroup_33_ready;
  wire       [21:0]   mulResGroup_33_payload;
  wire                mulResGroup_34_valid;
  wire                mulResGroup_34_ready;
  wire       [21:0]   mulResGroup_34_payload;
  wire                mulResGroup_35_valid;
  wire                mulResGroup_35_ready;
  wire       [21:0]   mulResGroup_35_payload;
  wire                mulResGroup_36_valid;
  wire                mulResGroup_36_ready;
  wire       [21:0]   mulResGroup_36_payload;
  wire                mulResGroup_37_valid;
  wire                mulResGroup_37_ready;
  wire       [21:0]   mulResGroup_37_payload;
  wire                mulResGroup_38_valid;
  wire                mulResGroup_38_ready;
  wire       [21:0]   mulResGroup_38_payload;
  wire                mulResGroup_39_valid;
  wire                mulResGroup_39_ready;
  wire       [21:0]   mulResGroup_39_payload;
  wire                mulResGroup_40_valid;
  wire                mulResGroup_40_ready;
  wire       [21:0]   mulResGroup_40_payload;
  wire                mulResGroup_41_valid;
  wire                mulResGroup_41_ready;
  wire       [21:0]   mulResGroup_41_payload;
  wire                mulResGroup_42_valid;
  wire                mulResGroup_42_ready;
  wire       [21:0]   mulResGroup_42_payload;
  wire                mulResGroup_43_valid;
  wire                mulResGroup_43_ready;
  wire       [21:0]   mulResGroup_43_payload;
  wire                mulResGroup_44_valid;
  wire                mulResGroup_44_ready;
  wire       [21:0]   mulResGroup_44_payload;
  wire                mulResGroup_45_valid;
  wire                mulResGroup_45_ready;
  wire       [21:0]   mulResGroup_45_payload;
  wire                mulResGroup_46_valid;
  wire                mulResGroup_46_ready;
  wire       [21:0]   mulResGroup_46_payload;
  wire                mulResGroup_47_valid;
  wire                mulResGroup_47_ready;
  wire       [21:0]   mulResGroup_47_payload;
  wire                mulResGroup_48_valid;
  wire                mulResGroup_48_ready;
  wire       [21:0]   mulResGroup_48_payload;
  wire                mulResGroup_49_valid;
  wire                mulResGroup_49_ready;
  wire       [21:0]   mulResGroup_49_payload;
  wire                mulResGroup_50_valid;
  wire                mulResGroup_50_ready;
  wire       [21:0]   mulResGroup_50_payload;
  wire                mulResGroup_51_valid;
  wire                mulResGroup_51_ready;
  wire       [21:0]   mulResGroup_51_payload;
  wire                mulResGroup_52_valid;
  wire                mulResGroup_52_ready;
  wire       [21:0]   mulResGroup_52_payload;
  wire                mulResGroup_53_valid;
  wire                mulResGroup_53_ready;
  wire       [21:0]   mulResGroup_53_payload;
  wire                mulResGroup_54_valid;
  wire                mulResGroup_54_ready;
  wire       [21:0]   mulResGroup_54_payload;
  wire                mulResGroup_55_valid;
  wire                mulResGroup_55_ready;
  wire       [21:0]   mulResGroup_55_payload;
  wire                mulResGroup_56_valid;
  wire                mulResGroup_56_ready;
  wire       [21:0]   mulResGroup_56_payload;
  wire                mulResGroup_57_valid;
  wire                mulResGroup_57_ready;
  wire       [21:0]   mulResGroup_57_payload;
  wire                mulResGroup_58_valid;
  wire                mulResGroup_58_ready;
  wire       [21:0]   mulResGroup_58_payload;
  wire                mulResGroup_59_valid;
  wire                mulResGroup_59_ready;
  wire       [21:0]   mulResGroup_59_payload;
  wire                mulResGroup_60_valid;
  wire                mulResGroup_60_ready;
  wire       [21:0]   mulResGroup_60_payload;
  wire                mulResGroup_61_valid;
  wire                mulResGroup_61_ready;
  wire       [21:0]   mulResGroup_61_payload;
  wire                mulResGroup_62_valid;
  wire                mulResGroup_62_ready;
  wire       [21:0]   mulResGroup_62_payload;
  wire                mulResGroup_63_valid;
  wire                mulResGroup_63_ready;
  wire       [21:0]   mulResGroup_63_payload;
  wire                mulResVec_valid;
  wire                mulResVec_ready;
  wire       [21:0]   mulResVec_payload_0;
  wire       [21:0]   mulResVec_payload_1;
  wire       [21:0]   mulResVec_payload_2;
  wire       [21:0]   mulResVec_payload_3;
  wire       [21:0]   mulResVec_payload_4;
  wire       [21:0]   mulResVec_payload_5;
  wire       [21:0]   mulResVec_payload_6;
  wire       [21:0]   mulResVec_payload_7;
  wire       [21:0]   mulResVec_payload_8;
  wire       [21:0]   mulResVec_payload_9;
  wire       [21:0]   mulResVec_payload_10;
  wire       [21:0]   mulResVec_payload_11;
  wire       [21:0]   mulResVec_payload_12;
  wire       [21:0]   mulResVec_payload_13;
  wire       [21:0]   mulResVec_payload_14;
  wire       [21:0]   mulResVec_payload_15;
  wire       [21:0]   mulResVec_payload_16;
  wire       [21:0]   mulResVec_payload_17;
  wire       [21:0]   mulResVec_payload_18;
  wire       [21:0]   mulResVec_payload_19;
  wire       [21:0]   mulResVec_payload_20;
  wire       [21:0]   mulResVec_payload_21;
  wire       [21:0]   mulResVec_payload_22;
  wire       [21:0]   mulResVec_payload_23;
  wire       [21:0]   mulResVec_payload_24;
  wire       [21:0]   mulResVec_payload_25;
  wire       [21:0]   mulResVec_payload_26;
  wire       [21:0]   mulResVec_payload_27;
  wire       [21:0]   mulResVec_payload_28;
  wire       [21:0]   mulResVec_payload_29;
  wire       [21:0]   mulResVec_payload_30;
  wire       [21:0]   mulResVec_payload_31;
  wire       [21:0]   mulResVec_payload_32;
  wire       [21:0]   mulResVec_payload_33;
  wire       [21:0]   mulResVec_payload_34;
  wire       [21:0]   mulResVec_payload_35;
  wire       [21:0]   mulResVec_payload_36;
  wire       [21:0]   mulResVec_payload_37;
  wire       [21:0]   mulResVec_payload_38;
  wire       [21:0]   mulResVec_payload_39;
  wire       [21:0]   mulResVec_payload_40;
  wire       [21:0]   mulResVec_payload_41;
  wire       [21:0]   mulResVec_payload_42;
  wire       [21:0]   mulResVec_payload_43;
  wire       [21:0]   mulResVec_payload_44;
  wire       [21:0]   mulResVec_payload_45;
  wire       [21:0]   mulResVec_payload_46;
  wire       [21:0]   mulResVec_payload_47;
  wire       [21:0]   mulResVec_payload_48;
  wire       [21:0]   mulResVec_payload_49;
  wire       [21:0]   mulResVec_payload_50;
  wire       [21:0]   mulResVec_payload_51;
  wire       [21:0]   mulResVec_payload_52;
  wire       [21:0]   mulResVec_payload_53;
  wire       [21:0]   mulResVec_payload_54;
  wire       [21:0]   mulResVec_payload_55;
  wire       [21:0]   mulResVec_payload_56;
  wire       [21:0]   mulResVec_payload_57;
  wire       [21:0]   mulResVec_payload_58;
  wire       [21:0]   mulResVec_payload_59;
  wire       [21:0]   mulResVec_payload_60;
  wire       [21:0]   mulResVec_payload_61;
  wire       [21:0]   mulResVec_payload_62;
  wire       [21:0]   mulResVec_payload_63;
  wire                mulResVec_translated_valid;
  wire                mulResVec_translated_ready;
  wire       [21:0]   mulResVec_translated_payload;

  assign _zz_mulResGroup_0_payload = 9'h0;
  assign _zz_mulResGroup_1_payload = 9'h0;
  assign _zz_mulResGroup_2_payload = 9'h0;
  assign _zz_mulResGroup_3_payload = 9'h0;
  assign _zz_mulResGroup_4_payload = 9'h0;
  assign _zz_mulResGroup_5_payload = 9'h0;
  assign _zz_mulResGroup_6_payload = 9'h0;
  assign _zz_mulResGroup_7_payload = 9'h0;
  assign _zz_mulResGroup_8_payload = 9'h0;
  assign _zz_mulResGroup_9_payload = 9'h0;
  assign _zz_mulResGroup_10_payload = 9'h0;
  assign _zz_mulResGroup_11_payload = 9'h0;
  assign _zz_mulResGroup_12_payload = 9'h0;
  assign _zz_mulResGroup_13_payload = 9'h0;
  assign _zz_mulResGroup_14_payload = 9'h0;
  assign _zz_mulResGroup_15_payload = 9'h0;
  assign _zz_mulResGroup_16_payload = ($signed(_zz_mulResGroup_16_payload_1) * $signed(_zz_mulResGroup_16_payload_2));
  assign _zz_mulResGroup_16_payload_1 = 1'b1;
  assign _zz_mulResGroup_16_payload_2 = ($signed(_zz_mulResGroup_16_payload_3) + $signed(_zz_mulResGroup_16_payload_4));
  assign _zz_mulResGroup_16_payload_3 = {{1{inputAll_16_fork_io_outputs_0_payload[7]}}, inputAll_16_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_16_payload_4 = {{1{inputAll_111_fork_io_outputs_0_payload[7]}}, inputAll_111_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_17_payload = ($signed(_zz_mulResGroup_17_payload_1) * $signed(_zz_mulResGroup_17_payload_2));
  assign _zz_mulResGroup_17_payload_1 = 1'b1;
  assign _zz_mulResGroup_17_payload_2 = ($signed(_zz_mulResGroup_17_payload_3) + $signed(_zz_mulResGroup_17_payload_4));
  assign _zz_mulResGroup_17_payload_3 = {{1{inputAll_17_fork_io_outputs_0_payload[7]}}, inputAll_17_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_17_payload_4 = {{1{inputAll_110_fork_io_outputs_0_payload[7]}}, inputAll_110_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_18_payload = ($signed(_zz_mulResGroup_18_payload_1) * $signed(_zz_mulResGroup_18_payload_2));
  assign _zz_mulResGroup_18_payload_1 = 1'b1;
  assign _zz_mulResGroup_18_payload_2 = ($signed(_zz_mulResGroup_18_payload_3) + $signed(_zz_mulResGroup_18_payload_4));
  assign _zz_mulResGroup_18_payload_3 = {{1{inputAll_18_fork_io_outputs_0_payload[7]}}, inputAll_18_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_18_payload_4 = {{1{inputAll_109_fork_io_outputs_0_payload[7]}}, inputAll_109_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_19_payload = 9'h0;
  assign _zz_mulResGroup_20_payload = 9'h0;
  assign _zz_mulResGroup_21_payload = ($signed(_zz_mulResGroup_21_payload_1) * $signed(_zz_mulResGroup_21_payload_2));
  assign _zz_mulResGroup_21_payload_1 = 2'b01;
  assign _zz_mulResGroup_21_payload_2 = ($signed(_zz_mulResGroup_21_payload_3) + $signed(_zz_mulResGroup_21_payload_4));
  assign _zz_mulResGroup_21_payload_3 = {{1{inputAll_21_fork_io_outputs_0_payload[7]}}, inputAll_21_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_21_payload_4 = {{1{inputAll_106_fork_io_outputs_0_payload[7]}}, inputAll_106_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_22_payload = ($signed(_zz_mulResGroup_22_payload_1) * $signed(_zz_mulResGroup_22_payload_2));
  assign _zz_mulResGroup_22_payload_1 = 2'b01;
  assign _zz_mulResGroup_22_payload_2 = ($signed(_zz_mulResGroup_22_payload_3) + $signed(_zz_mulResGroup_22_payload_4));
  assign _zz_mulResGroup_22_payload_3 = {{1{inputAll_22_fork_io_outputs_0_payload[7]}}, inputAll_22_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_22_payload_4 = {{1{inputAll_105_fork_io_outputs_0_payload[7]}}, inputAll_105_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_23_payload = ($signed(_zz_mulResGroup_23_payload_1) * $signed(_zz_mulResGroup_23_payload_2));
  assign _zz_mulResGroup_23_payload_1 = 2'b01;
  assign _zz_mulResGroup_23_payload_2 = ($signed(_zz_mulResGroup_23_payload_3) + $signed(_zz_mulResGroup_23_payload_4));
  assign _zz_mulResGroup_23_payload_3 = {{1{inputAll_23_fork_io_outputs_0_payload[7]}}, inputAll_23_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_23_payload_4 = {{1{inputAll_104_fork_io_outputs_0_payload[7]}}, inputAll_104_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_24_payload = ($signed(_zz_mulResGroup_24_payload_1) * $signed(_zz_mulResGroup_24_payload_2));
  assign _zz_mulResGroup_24_payload_1 = 2'b01;
  assign _zz_mulResGroup_24_payload_2 = ($signed(_zz_mulResGroup_24_payload_3) + $signed(_zz_mulResGroup_24_payload_4));
  assign _zz_mulResGroup_24_payload_3 = {{1{inputAll_24_fork_io_outputs_0_payload[7]}}, inputAll_24_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_24_payload_4 = {{1{inputAll_103_fork_io_outputs_0_payload[7]}}, inputAll_103_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_25_payload = ($signed(_zz_mulResGroup_25_payload_1) * $signed(_zz_mulResGroup_25_payload_2));
  assign _zz_mulResGroup_25_payload_1 = 2'b01;
  assign _zz_mulResGroup_25_payload_2 = ($signed(_zz_mulResGroup_25_payload_3) + $signed(_zz_mulResGroup_25_payload_4));
  assign _zz_mulResGroup_25_payload_3 = {{1{inputAll_25_fork_io_outputs_0_payload[7]}}, inputAll_25_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_25_payload_4 = {{1{inputAll_102_fork_io_outputs_0_payload[7]}}, inputAll_102_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_26_payload = 9'h0;
  assign _zz_mulResGroup_27_payload = ($signed(_zz_mulResGroup_27_payload_1) * $signed(_zz_mulResGroup_27_payload_2));
  assign _zz_mulResGroup_27_payload_1 = 1'b1;
  assign _zz_mulResGroup_27_payload_2 = ($signed(_zz_mulResGroup_27_payload_3) + $signed(_zz_mulResGroup_27_payload_4));
  assign _zz_mulResGroup_27_payload_3 = {{1{inputAll_27_fork_io_outputs_0_payload[7]}}, inputAll_27_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_27_payload_4 = {{1{inputAll_100_fork_io_outputs_0_payload[7]}}, inputAll_100_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_28_payload = ($signed(_zz_mulResGroup_28_payload_1) * $signed(_zz_mulResGroup_28_payload_2));
  assign _zz_mulResGroup_28_payload_1 = 2'b10;
  assign _zz_mulResGroup_28_payload_2 = ($signed(_zz_mulResGroup_28_payload_3) + $signed(_zz_mulResGroup_28_payload_4));
  assign _zz_mulResGroup_28_payload_3 = {{1{inputAll_28_fork_io_outputs_0_payload[7]}}, inputAll_28_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_28_payload_4 = {{1{inputAll_99_fork_io_outputs_0_payload[7]}}, inputAll_99_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_29_payload = ($signed(_zz_mulResGroup_29_payload_1) * $signed(_zz_mulResGroup_29_payload_2));
  assign _zz_mulResGroup_29_payload_1 = 2'b10;
  assign _zz_mulResGroup_29_payload_2 = ($signed(_zz_mulResGroup_29_payload_3) + $signed(_zz_mulResGroup_29_payload_4));
  assign _zz_mulResGroup_29_payload_3 = {{1{inputAll_29_fork_io_outputs_0_payload[7]}}, inputAll_29_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_29_payload_4 = {{1{inputAll_98_fork_io_outputs_0_payload[7]}}, inputAll_98_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_30_payload = ($signed(_zz_mulResGroup_30_payload_1) * $signed(_zz_mulResGroup_30_payload_2));
  assign _zz_mulResGroup_30_payload_1 = 2'b10;
  assign _zz_mulResGroup_30_payload_2 = ($signed(_zz_mulResGroup_30_payload_3) + $signed(_zz_mulResGroup_30_payload_4));
  assign _zz_mulResGroup_30_payload_3 = {{1{inputAll_30_fork_io_outputs_0_payload[7]}}, inputAll_30_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_30_payload_4 = {{1{inputAll_97_fork_io_outputs_0_payload[7]}}, inputAll_97_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_31_payload = ($signed(_zz_mulResGroup_31_payload_1) * $signed(_zz_mulResGroup_31_payload_2));
  assign _zz_mulResGroup_31_payload_1 = 2'b10;
  assign _zz_mulResGroup_31_payload_2 = ($signed(_zz_mulResGroup_31_payload_3) + $signed(_zz_mulResGroup_31_payload_4));
  assign _zz_mulResGroup_31_payload_3 = {{1{inputAll_31_fork_io_outputs_0_payload[7]}}, inputAll_31_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_31_payload_4 = {{1{inputAll_96_fork_io_outputs_0_payload[7]}}, inputAll_96_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_32_payload = 9'h0;
  assign _zz_mulResGroup_33_payload = ($signed(_zz_mulResGroup_33_payload_1) * $signed(_zz_mulResGroup_33_payload_2));
  assign _zz_mulResGroup_33_payload_1 = 2'b01;
  assign _zz_mulResGroup_33_payload_2 = ($signed(_zz_mulResGroup_33_payload_3) + $signed(_zz_mulResGroup_33_payload_4));
  assign _zz_mulResGroup_33_payload_3 = {{1{inputAll_33_fork_io_outputs_0_payload[7]}}, inputAll_33_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_33_payload_4 = {{1{inputAll_94_fork_io_outputs_0_payload[7]}}, inputAll_94_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_34_payload = ($signed(_zz_mulResGroup_34_payload_1) * $signed(_zz_mulResGroup_34_payload_2));
  assign _zz_mulResGroup_34_payload_1 = 3'b011;
  assign _zz_mulResGroup_34_payload_2 = ($signed(_zz_mulResGroup_34_payload_3) + $signed(_zz_mulResGroup_34_payload_4));
  assign _zz_mulResGroup_34_payload_3 = {{1{inputAll_34_fork_io_outputs_0_payload[7]}}, inputAll_34_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_34_payload_4 = {{1{inputAll_93_fork_io_outputs_0_payload[7]}}, inputAll_93_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_35_payload = ($signed(_zz_mulResGroup_35_payload_1) * $signed(_zz_mulResGroup_35_payload_2));
  assign _zz_mulResGroup_35_payload_1 = 3'b011;
  assign _zz_mulResGroup_35_payload_2 = ($signed(_zz_mulResGroup_35_payload_3) + $signed(_zz_mulResGroup_35_payload_4));
  assign _zz_mulResGroup_35_payload_3 = {{1{inputAll_35_fork_io_outputs_0_payload[7]}}, inputAll_35_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_35_payload_4 = {{1{inputAll_92_fork_io_outputs_0_payload[7]}}, inputAll_92_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_36_payload = ($signed(_zz_mulResGroup_36_payload_1) * $signed(_zz_mulResGroup_36_payload_2));
  assign _zz_mulResGroup_36_payload_1 = 4'b0100;
  assign _zz_mulResGroup_36_payload_2 = ($signed(_zz_mulResGroup_36_payload_3) + $signed(_zz_mulResGroup_36_payload_4));
  assign _zz_mulResGroup_36_payload_3 = {{1{inputAll_36_fork_io_outputs_0_payload[7]}}, inputAll_36_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_36_payload_4 = {{1{inputAll_91_fork_io_outputs_0_payload[7]}}, inputAll_91_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_37_payload = ($signed(_zz_mulResGroup_37_payload_1) * $signed(_zz_mulResGroup_37_payload_2));
  assign _zz_mulResGroup_37_payload_1 = 3'b011;
  assign _zz_mulResGroup_37_payload_2 = ($signed(_zz_mulResGroup_37_payload_3) + $signed(_zz_mulResGroup_37_payload_4));
  assign _zz_mulResGroup_37_payload_3 = {{1{inputAll_37_fork_io_outputs_0_payload[7]}}, inputAll_37_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_37_payload_4 = {{1{inputAll_90_fork_io_outputs_0_payload[7]}}, inputAll_90_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_38_payload = ($signed(_zz_mulResGroup_38_payload_1) * $signed(_zz_mulResGroup_38_payload_2));
  assign _zz_mulResGroup_38_payload_1 = 2'b01;
  assign _zz_mulResGroup_38_payload_2 = ($signed(_zz_mulResGroup_38_payload_3) + $signed(_zz_mulResGroup_38_payload_4));
  assign _zz_mulResGroup_38_payload_3 = {{1{inputAll_38_fork_io_outputs_0_payload[7]}}, inputAll_38_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_38_payload_4 = {{1{inputAll_89_fork_io_outputs_0_payload[7]}}, inputAll_89_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_39_payload = ($signed(_zz_mulResGroup_39_payload_1) * $signed(_zz_mulResGroup_39_payload_2));
  assign _zz_mulResGroup_39_payload_1 = 1'b1;
  assign _zz_mulResGroup_39_payload_2 = ($signed(_zz_mulResGroup_39_payload_3) + $signed(_zz_mulResGroup_39_payload_4));
  assign _zz_mulResGroup_39_payload_3 = {{1{inputAll_39_fork_io_outputs_0_payload[7]}}, inputAll_39_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_39_payload_4 = {{1{inputAll_88_fork_io_outputs_0_payload[7]}}, inputAll_88_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_40_payload = ($signed(_zz_mulResGroup_40_payload_1) * $signed(_zz_mulResGroup_40_payload_2));
  assign _zz_mulResGroup_40_payload_1 = 3'b101;
  assign _zz_mulResGroup_40_payload_2 = ($signed(_zz_mulResGroup_40_payload_3) + $signed(_zz_mulResGroup_40_payload_4));
  assign _zz_mulResGroup_40_payload_3 = {{1{inputAll_40_fork_io_outputs_0_payload[7]}}, inputAll_40_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_40_payload_4 = {{1{inputAll_87_fork_io_outputs_0_payload[7]}}, inputAll_87_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_41_payload = ($signed(_zz_mulResGroup_41_payload_1) * $signed(_zz_mulResGroup_41_payload_2));
  assign _zz_mulResGroup_41_payload_1 = 4'b1011;
  assign _zz_mulResGroup_41_payload_2 = ($signed(_zz_mulResGroup_41_payload_3) + $signed(_zz_mulResGroup_41_payload_4));
  assign _zz_mulResGroup_41_payload_3 = {{1{inputAll_41_fork_io_outputs_0_payload[7]}}, inputAll_41_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_41_payload_4 = {{1{inputAll_86_fork_io_outputs_0_payload[7]}}, inputAll_86_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_42_payload = ($signed(_zz_mulResGroup_42_payload_1) * $signed(_zz_mulResGroup_42_payload_2));
  assign _zz_mulResGroup_42_payload_1 = 4'b1010;
  assign _zz_mulResGroup_42_payload_2 = ($signed(_zz_mulResGroup_42_payload_3) + $signed(_zz_mulResGroup_42_payload_4));
  assign _zz_mulResGroup_42_payload_3 = {{1{inputAll_42_fork_io_outputs_0_payload[7]}}, inputAll_42_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_42_payload_4 = {{1{inputAll_85_fork_io_outputs_0_payload[7]}}, inputAll_85_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_43_payload = ($signed(_zz_mulResGroup_43_payload_1) * $signed(_zz_mulResGroup_43_payload_2));
  assign _zz_mulResGroup_43_payload_1 = 4'b1011;
  assign _zz_mulResGroup_43_payload_2 = ($signed(_zz_mulResGroup_43_payload_3) + $signed(_zz_mulResGroup_43_payload_4));
  assign _zz_mulResGroup_43_payload_3 = {{1{inputAll_43_fork_io_outputs_0_payload[7]}}, inputAll_43_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_43_payload_4 = {{1{inputAll_84_fork_io_outputs_0_payload[7]}}, inputAll_84_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_44_payload = ($signed(_zz_mulResGroup_44_payload_1) * $signed(_zz_mulResGroup_44_payload_2));
  assign _zz_mulResGroup_44_payload_1 = 2'b10;
  assign _zz_mulResGroup_44_payload_2 = ($signed(_zz_mulResGroup_44_payload_3) + $signed(_zz_mulResGroup_44_payload_4));
  assign _zz_mulResGroup_44_payload_3 = {{1{inputAll_44_fork_io_outputs_0_payload[7]}}, inputAll_44_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_44_payload_4 = {{1{inputAll_83_fork_io_outputs_0_payload[7]}}, inputAll_83_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_45_payload = ($signed(_zz_mulResGroup_45_payload_1) * $signed(_zz_mulResGroup_45_payload_2));
  assign _zz_mulResGroup_45_payload_1 = 2'b01;
  assign _zz_mulResGroup_45_payload_2 = ($signed(_zz_mulResGroup_45_payload_3) + $signed(_zz_mulResGroup_45_payload_4));
  assign _zz_mulResGroup_45_payload_3 = {{1{inputAll_45_fork_io_outputs_0_payload[7]}}, inputAll_45_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_45_payload_4 = {{1{inputAll_82_fork_io_outputs_0_payload[7]}}, inputAll_82_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_46_payload = ($signed(_zz_mulResGroup_46_payload_1) * $signed(_zz_mulResGroup_46_payload_2));
  assign _zz_mulResGroup_46_payload_1 = 4'b0101;
  assign _zz_mulResGroup_46_payload_2 = ($signed(_zz_mulResGroup_46_payload_3) + $signed(_zz_mulResGroup_46_payload_4));
  assign _zz_mulResGroup_46_payload_3 = {{1{inputAll_46_fork_io_outputs_0_payload[7]}}, inputAll_46_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_46_payload_4 = {{1{inputAll_81_fork_io_outputs_0_payload[7]}}, inputAll_81_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_47_payload = ($signed(_zz_mulResGroup_47_payload_1) * $signed(_zz_mulResGroup_47_payload_2));
  assign _zz_mulResGroup_47_payload_1 = 5'h08;
  assign _zz_mulResGroup_47_payload_2 = ($signed(_zz_mulResGroup_47_payload_3) + $signed(_zz_mulResGroup_47_payload_4));
  assign _zz_mulResGroup_47_payload_3 = {{1{inputAll_47_fork_io_outputs_0_payload[7]}}, inputAll_47_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_47_payload_4 = {{1{inputAll_80_fork_io_outputs_0_payload[7]}}, inputAll_80_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_48_payload = ($signed(_zz_mulResGroup_48_payload_1) * $signed(_zz_mulResGroup_48_payload_2));
  assign _zz_mulResGroup_48_payload_1 = 5'h09;
  assign _zz_mulResGroup_48_payload_2 = ($signed(_zz_mulResGroup_48_payload_3) + $signed(_zz_mulResGroup_48_payload_4));
  assign _zz_mulResGroup_48_payload_3 = {{1{inputAll_48_fork_io_outputs_0_payload[7]}}, inputAll_48_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_48_payload_4 = {{1{inputAll_79_fork_io_outputs_0_payload[7]}}, inputAll_79_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_49_payload = ($signed(_zz_mulResGroup_49_payload_1) * $signed(_zz_mulResGroup_49_payload_2));
  assign _zz_mulResGroup_49_payload_1 = 5'h08;
  assign _zz_mulResGroup_49_payload_2 = ($signed(_zz_mulResGroup_49_payload_3) + $signed(_zz_mulResGroup_49_payload_4));
  assign _zz_mulResGroup_49_payload_3 = {{1{inputAll_49_fork_io_outputs_0_payload[7]}}, inputAll_49_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_49_payload_4 = {{1{inputAll_78_fork_io_outputs_0_payload[7]}}, inputAll_78_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_50_payload = ($signed(_zz_mulResGroup_50_payload_1) * $signed(_zz_mulResGroup_50_payload_2));
  assign _zz_mulResGroup_50_payload_1 = 4'b0101;
  assign _zz_mulResGroup_50_payload_2 = ($signed(_zz_mulResGroup_50_payload_3) + $signed(_zz_mulResGroup_50_payload_4));
  assign _zz_mulResGroup_50_payload_3 = {{1{inputAll_50_fork_io_outputs_0_payload[7]}}, inputAll_50_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_50_payload_4 = {{1{inputAll_77_fork_io_outputs_0_payload[7]}}, inputAll_77_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_51_payload = 9'h0;
  assign _zz_mulResGroup_52_payload = ($signed(_zz_mulResGroup_52_payload_1) * $signed(_zz_mulResGroup_52_payload_2));
  assign _zz_mulResGroup_52_payload_1 = 4'b1010;
  assign _zz_mulResGroup_52_payload_2 = ($signed(_zz_mulResGroup_52_payload_3) + $signed(_zz_mulResGroup_52_payload_4));
  assign _zz_mulResGroup_52_payload_3 = {{1{inputAll_52_fork_io_outputs_0_payload[7]}}, inputAll_52_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_52_payload_4 = {{1{inputAll_75_fork_io_outputs_0_payload[7]}}, inputAll_75_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_53_payload = ($signed(_zz_mulResGroup_53_payload_1) * $signed(_zz_mulResGroup_53_payload_2));
  assign _zz_mulResGroup_53_payload_1 = 5'h14;
  assign _zz_mulResGroup_53_payload_2 = ($signed(_zz_mulResGroup_53_payload_3) + $signed(_zz_mulResGroup_53_payload_4));
  assign _zz_mulResGroup_53_payload_3 = {{1{inputAll_53_fork_io_outputs_0_payload[7]}}, inputAll_53_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_53_payload_4 = {{1{inputAll_74_fork_io_outputs_0_payload[7]}}, inputAll_74_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_54_payload = ($signed(_zz_mulResGroup_54_payload_1) * $signed(_zz_mulResGroup_54_payload_2));
  assign _zz_mulResGroup_54_payload_1 = 5'h10;
  assign _zz_mulResGroup_54_payload_2 = ($signed(_zz_mulResGroup_54_payload_3) + $signed(_zz_mulResGroup_54_payload_4));
  assign _zz_mulResGroup_54_payload_3 = {{1{inputAll_54_fork_io_outputs_0_payload[7]}}, inputAll_54_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_54_payload_4 = {{1{inputAll_73_fork_io_outputs_0_payload[7]}}, inputAll_73_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_55_payload = ($signed(_zz_mulResGroup_55_payload_1) * $signed(_zz_mulResGroup_55_payload_2));
  assign _zz_mulResGroup_55_payload_1 = 6'h2f;
  assign _zz_mulResGroup_55_payload_2 = ($signed(_zz_mulResGroup_55_payload_3) + $signed(_zz_mulResGroup_55_payload_4));
  assign _zz_mulResGroup_55_payload_3 = {{1{inputAll_55_fork_io_outputs_0_payload[7]}}, inputAll_55_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_55_payload_4 = {{1{inputAll_72_fork_io_outputs_0_payload[7]}}, inputAll_72_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_56_payload = ($signed(_zz_mulResGroup_56_payload_1) * $signed(_zz_mulResGroup_56_payload_2));
  assign _zz_mulResGroup_56_payload_1 = 5'h14;
  assign _zz_mulResGroup_56_payload_2 = ($signed(_zz_mulResGroup_56_payload_3) + $signed(_zz_mulResGroup_56_payload_4));
  assign _zz_mulResGroup_56_payload_3 = {{1{inputAll_56_fork_io_outputs_0_payload[7]}}, inputAll_56_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_56_payload_4 = {{1{inputAll_71_fork_io_outputs_0_payload[7]}}, inputAll_71_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_57_payload = ($signed(_zz_mulResGroup_57_payload_1) * $signed(_zz_mulResGroup_57_payload_2));
  assign _zz_mulResGroup_57_payload_1 = 3'b101;
  assign _zz_mulResGroup_57_payload_2 = ($signed(_zz_mulResGroup_57_payload_3) + $signed(_zz_mulResGroup_57_payload_4));
  assign _zz_mulResGroup_57_payload_3 = {{1{inputAll_57_fork_io_outputs_0_payload[7]}}, inputAll_57_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_57_payload_4 = {{1{inputAll_70_fork_io_outputs_0_payload[7]}}, inputAll_70_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_58_payload = ($signed(_zz_mulResGroup_58_payload_1) * $signed(_zz_mulResGroup_58_payload_2));
  assign _zz_mulResGroup_58_payload_1 = 5'h0b;
  assign _zz_mulResGroup_58_payload_2 = ($signed(_zz_mulResGroup_58_payload_3) + $signed(_zz_mulResGroup_58_payload_4));
  assign _zz_mulResGroup_58_payload_3 = {{1{inputAll_58_fork_io_outputs_0_payload[7]}}, inputAll_58_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_58_payload_4 = {{1{inputAll_69_fork_io_outputs_0_payload[7]}}, inputAll_69_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_59_payload = ($signed(_zz_mulResGroup_59_payload_1) * $signed(_zz_mulResGroup_59_payload_2));
  assign _zz_mulResGroup_59_payload_1 = 6'h1c;
  assign _zz_mulResGroup_59_payload_2 = ($signed(_zz_mulResGroup_59_payload_3) + $signed(_zz_mulResGroup_59_payload_4));
  assign _zz_mulResGroup_59_payload_3 = {{1{inputAll_59_fork_io_outputs_0_payload[7]}}, inputAll_59_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_59_payload_4 = {{1{inputAll_68_fork_io_outputs_0_payload[7]}}, inputAll_68_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_60_payload = ($signed(_zz_mulResGroup_60_payload_1) * $signed(_zz_mulResGroup_60_payload_2));
  assign _zz_mulResGroup_60_payload_1 = 7'h2d;
  assign _zz_mulResGroup_60_payload_2 = ($signed(_zz_mulResGroup_60_payload_3) + $signed(_zz_mulResGroup_60_payload_4));
  assign _zz_mulResGroup_60_payload_3 = {{1{inputAll_60_fork_io_outputs_0_payload[7]}}, inputAll_60_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_60_payload_4 = {{1{inputAll_67_fork_io_outputs_0_payload[7]}}, inputAll_67_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_61_payload = ($signed(_zz_mulResGroup_61_payload_1) * $signed(_zz_mulResGroup_61_payload_2));
  assign _zz_mulResGroup_61_payload_1 = 7'h3e;
  assign _zz_mulResGroup_61_payload_2 = ($signed(_zz_mulResGroup_61_payload_3) + $signed(_zz_mulResGroup_61_payload_4));
  assign _zz_mulResGroup_61_payload_3 = {{1{inputAll_61_fork_io_outputs_0_payload[7]}}, inputAll_61_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_61_payload_4 = {{1{inputAll_66_fork_io_outputs_0_payload[7]}}, inputAll_66_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_62_payload = ($signed(_zz_mulResGroup_62_payload_1) * $signed(_zz_mulResGroup_62_payload_2));
  assign _zz_mulResGroup_62_payload_1 = 8'h4a;
  assign _zz_mulResGroup_62_payload_2 = ($signed(_zz_mulResGroup_62_payload_3) + $signed(_zz_mulResGroup_62_payload_4));
  assign _zz_mulResGroup_62_payload_3 = {{1{inputAll_62_fork_io_outputs_0_payload[7]}}, inputAll_62_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_62_payload_4 = {{1{inputAll_65_fork_io_outputs_0_payload[7]}}, inputAll_65_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_63_payload = ($signed(_zz_mulResGroup_63_payload_1) * $signed(_zz_mulResGroup_63_payload_2));
  assign _zz_mulResGroup_63_payload_1 = 8'h51;
  assign _zz_mulResGroup_63_payload_2 = ($signed(_zz_mulResGroup_63_payload_3) + $signed(_zz_mulResGroup_63_payload_4));
  assign _zz_mulResGroup_63_payload_3 = {{1{inputAll_63_fork_io_outputs_0_payload[7]}}, inputAll_63_fork_io_outputs_0_payload};
  assign _zz_mulResGroup_63_payload_4 = {{1{inputAll_64_fork_io_outputs_0_payload[7]}}, inputAll_64_fork_io_outputs_0_payload};
  assign _zz_mulResVec_translated_payload = ($signed(_zz_mulResVec_translated_payload_1) + $signed(_zz_mulResVec_translated_payload_16));
  assign _zz_mulResVec_translated_payload_1 = ($signed(_zz_mulResVec_translated_payload_2) + $signed(_zz_mulResVec_translated_payload_9));
  assign _zz_mulResVec_translated_payload_2 = ($signed(_zz_mulResVec_translated_payload_3) + $signed(_zz_mulResVec_translated_payload_6));
  assign _zz_mulResVec_translated_payload_3 = ($signed(_zz_mulResVec_translated_payload_4) + $signed(_zz_mulResVec_translated_payload_5));
  assign _zz_mulResVec_translated_payload_4 = ($signed(mulResVec_payload_0) + $signed(mulResVec_payload_1));
  assign _zz_mulResVec_translated_payload_5 = ($signed(mulResVec_payload_2) + $signed(mulResVec_payload_3));
  assign _zz_mulResVec_translated_payload_6 = ($signed(_zz_mulResVec_translated_payload_7) + $signed(_zz_mulResVec_translated_payload_8));
  assign _zz_mulResVec_translated_payload_7 = ($signed(mulResVec_payload_4) + $signed(mulResVec_payload_5));
  assign _zz_mulResVec_translated_payload_8 = ($signed(mulResVec_payload_6) + $signed(mulResVec_payload_7));
  assign _zz_mulResVec_translated_payload_9 = ($signed(_zz_mulResVec_translated_payload_10) + $signed(_zz_mulResVec_translated_payload_13));
  assign _zz_mulResVec_translated_payload_10 = ($signed(_zz_mulResVec_translated_payload_11) + $signed(_zz_mulResVec_translated_payload_12));
  assign _zz_mulResVec_translated_payload_11 = ($signed(mulResVec_payload_8) + $signed(mulResVec_payload_9));
  assign _zz_mulResVec_translated_payload_12 = ($signed(mulResVec_payload_10) + $signed(mulResVec_payload_11));
  assign _zz_mulResVec_translated_payload_13 = ($signed(_zz_mulResVec_translated_payload_14) + $signed(_zz_mulResVec_translated_payload_15));
  assign _zz_mulResVec_translated_payload_14 = ($signed(mulResVec_payload_12) + $signed(mulResVec_payload_13));
  assign _zz_mulResVec_translated_payload_15 = ($signed(mulResVec_payload_14) + $signed(mulResVec_payload_15));
  assign _zz_mulResVec_translated_payload_16 = ($signed(_zz_mulResVec_translated_payload_17) + $signed(_zz_mulResVec_translated_payload_24));
  assign _zz_mulResVec_translated_payload_17 = ($signed(_zz_mulResVec_translated_payload_18) + $signed(_zz_mulResVec_translated_payload_21));
  assign _zz_mulResVec_translated_payload_18 = ($signed(_zz_mulResVec_translated_payload_19) + $signed(_zz_mulResVec_translated_payload_20));
  assign _zz_mulResVec_translated_payload_19 = ($signed(mulResVec_payload_16) + $signed(mulResVec_payload_17));
  assign _zz_mulResVec_translated_payload_20 = ($signed(mulResVec_payload_18) + $signed(mulResVec_payload_19));
  assign _zz_mulResVec_translated_payload_21 = ($signed(_zz_mulResVec_translated_payload_22) + $signed(_zz_mulResVec_translated_payload_23));
  assign _zz_mulResVec_translated_payload_22 = ($signed(mulResVec_payload_20) + $signed(mulResVec_payload_21));
  assign _zz_mulResVec_translated_payload_23 = ($signed(mulResVec_payload_22) + $signed(mulResVec_payload_23));
  assign _zz_mulResVec_translated_payload_24 = ($signed(_zz_mulResVec_translated_payload_25) + $signed(_zz_mulResVec_translated_payload_28));
  assign _zz_mulResVec_translated_payload_25 = ($signed(_zz_mulResVec_translated_payload_26) + $signed(_zz_mulResVec_translated_payload_27));
  assign _zz_mulResVec_translated_payload_26 = ($signed(mulResVec_payload_24) + $signed(mulResVec_payload_25));
  assign _zz_mulResVec_translated_payload_27 = ($signed(mulResVec_payload_26) + $signed(mulResVec_payload_27));
  assign _zz_mulResVec_translated_payload_28 = ($signed(_zz_mulResVec_translated_payload_29) + $signed(_zz_mulResVec_translated_payload_30));
  assign _zz_mulResVec_translated_payload_29 = ($signed(mulResVec_payload_28) + $signed(mulResVec_payload_29));
  assign _zz_mulResVec_translated_payload_30 = ($signed(mulResVec_payload_30) + $signed(mulResVec_payload_31));
  assign _zz_mulResVec_translated_payload_31 = ($signed(_zz_mulResVec_translated_payload_32) + $signed(_zz_mulResVec_translated_payload_47));
  assign _zz_mulResVec_translated_payload_32 = ($signed(_zz_mulResVec_translated_payload_33) + $signed(_zz_mulResVec_translated_payload_40));
  assign _zz_mulResVec_translated_payload_33 = ($signed(_zz_mulResVec_translated_payload_34) + $signed(_zz_mulResVec_translated_payload_37));
  assign _zz_mulResVec_translated_payload_34 = ($signed(_zz_mulResVec_translated_payload_35) + $signed(_zz_mulResVec_translated_payload_36));
  assign _zz_mulResVec_translated_payload_35 = ($signed(mulResVec_payload_32) + $signed(mulResVec_payload_33));
  assign _zz_mulResVec_translated_payload_36 = ($signed(mulResVec_payload_34) + $signed(mulResVec_payload_35));
  assign _zz_mulResVec_translated_payload_37 = ($signed(_zz_mulResVec_translated_payload_38) + $signed(_zz_mulResVec_translated_payload_39));
  assign _zz_mulResVec_translated_payload_38 = ($signed(mulResVec_payload_36) + $signed(mulResVec_payload_37));
  assign _zz_mulResVec_translated_payload_39 = ($signed(mulResVec_payload_38) + $signed(mulResVec_payload_39));
  assign _zz_mulResVec_translated_payload_40 = ($signed(_zz_mulResVec_translated_payload_41) + $signed(_zz_mulResVec_translated_payload_44));
  assign _zz_mulResVec_translated_payload_41 = ($signed(_zz_mulResVec_translated_payload_42) + $signed(_zz_mulResVec_translated_payload_43));
  assign _zz_mulResVec_translated_payload_42 = ($signed(mulResVec_payload_40) + $signed(mulResVec_payload_41));
  assign _zz_mulResVec_translated_payload_43 = ($signed(mulResVec_payload_42) + $signed(mulResVec_payload_43));
  assign _zz_mulResVec_translated_payload_44 = ($signed(_zz_mulResVec_translated_payload_45) + $signed(_zz_mulResVec_translated_payload_46));
  assign _zz_mulResVec_translated_payload_45 = ($signed(mulResVec_payload_44) + $signed(mulResVec_payload_45));
  assign _zz_mulResVec_translated_payload_46 = ($signed(mulResVec_payload_46) + $signed(mulResVec_payload_47));
  assign _zz_mulResVec_translated_payload_47 = ($signed(_zz_mulResVec_translated_payload_48) + $signed(_zz_mulResVec_translated_payload_55));
  assign _zz_mulResVec_translated_payload_48 = ($signed(_zz_mulResVec_translated_payload_49) + $signed(_zz_mulResVec_translated_payload_52));
  assign _zz_mulResVec_translated_payload_49 = ($signed(_zz_mulResVec_translated_payload_50) + $signed(_zz_mulResVec_translated_payload_51));
  assign _zz_mulResVec_translated_payload_50 = ($signed(mulResVec_payload_48) + $signed(mulResVec_payload_49));
  assign _zz_mulResVec_translated_payload_51 = ($signed(mulResVec_payload_50) + $signed(mulResVec_payload_51));
  assign _zz_mulResVec_translated_payload_52 = ($signed(_zz_mulResVec_translated_payload_53) + $signed(_zz_mulResVec_translated_payload_54));
  assign _zz_mulResVec_translated_payload_53 = ($signed(mulResVec_payload_52) + $signed(mulResVec_payload_53));
  assign _zz_mulResVec_translated_payload_54 = ($signed(mulResVec_payload_54) + $signed(mulResVec_payload_55));
  assign _zz_mulResVec_translated_payload_55 = ($signed(_zz_mulResVec_translated_payload_56) + $signed(_zz_mulResVec_translated_payload_59));
  assign _zz_mulResVec_translated_payload_56 = ($signed(_zz_mulResVec_translated_payload_57) + $signed(_zz_mulResVec_translated_payload_58));
  assign _zz_mulResVec_translated_payload_57 = ($signed(mulResVec_payload_56) + $signed(mulResVec_payload_57));
  assign _zz_mulResVec_translated_payload_58 = ($signed(mulResVec_payload_58) + $signed(mulResVec_payload_59));
  assign _zz_mulResVec_translated_payload_59 = ($signed(_zz_mulResVec_translated_payload_60) + $signed(_zz_mulResVec_translated_payload_61));
  assign _zz_mulResVec_translated_payload_60 = ($signed(mulResVec_payload_60) + $signed(mulResVec_payload_61));
  assign _zz_mulResVec_translated_payload_61 = ($signed(mulResVec_payload_62) + $signed(mulResVec_payload_63));
  assign _zz_mulResVec_valid = ((((((((((((((((_zz_mulResVec_valid_1 && mulResGroup_32_valid) && mulResGroup_33_valid) && mulResGroup_34_valid) && mulResGroup_35_valid) && mulResGroup_36_valid) && mulResGroup_37_valid) && mulResGroup_38_valid) && mulResGroup_39_valid) && mulResGroup_40_valid) && mulResGroup_41_valid) && mulResGroup_42_valid) && mulResGroup_43_valid) && mulResGroup_44_valid) && mulResGroup_45_valid) && mulResGroup_46_valid) && mulResGroup_47_valid);
  assign _zz_mulResVec_valid_1 = ((((((((((((((((_zz_mulResVec_valid_2 && mulResGroup_16_valid) && mulResGroup_17_valid) && mulResGroup_18_valid) && mulResGroup_19_valid) && mulResGroup_20_valid) && mulResGroup_21_valid) && mulResGroup_22_valid) && mulResGroup_23_valid) && mulResGroup_24_valid) && mulResGroup_25_valid) && mulResGroup_26_valid) && mulResGroup_27_valid) && mulResGroup_28_valid) && mulResGroup_29_valid) && mulResGroup_30_valid) && mulResGroup_31_valid);
  assign _zz_mulResVec_valid_2 = (((((((((((((((mulResGroup_0_valid && mulResGroup_1_valid) && mulResGroup_2_valid) && mulResGroup_3_valid) && mulResGroup_4_valid) && mulResGroup_5_valid) && mulResGroup_6_valid) && mulResGroup_7_valid) && mulResGroup_8_valid) && mulResGroup_9_valid) && mulResGroup_10_valid) && mulResGroup_11_valid) && mulResGroup_12_valid) && mulResGroup_13_valid) && mulResGroup_14_valid) && mulResGroup_15_valid);
  StreamFork inputAll_0_fork (
    .io_input_valid          (inputAll_0_valid                      ), //i
    .io_input_ready          (inputAll_0_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_0_payload                    ), //i
    .io_outputs_0_valid      (inputAll_0_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_0_ready                   ), //i
    .io_outputs_0_payload    (inputAll_0_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_0_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_0_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_0_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_1_fork (
    .io_input_valid          (inputAll_1_valid                      ), //i
    .io_input_ready          (inputAll_1_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_1_payload                    ), //i
    .io_outputs_0_valid      (inputAll_1_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_1_ready                   ), //i
    .io_outputs_0_payload    (inputAll_1_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_1_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_1_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_1_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_2_fork (
    .io_input_valid          (inputAll_2_valid                      ), //i
    .io_input_ready          (inputAll_2_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_2_payload                    ), //i
    .io_outputs_0_valid      (inputAll_2_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_2_ready                   ), //i
    .io_outputs_0_payload    (inputAll_2_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_2_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_2_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_2_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_3_fork (
    .io_input_valid          (inputAll_3_valid                      ), //i
    .io_input_ready          (inputAll_3_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_3_payload                    ), //i
    .io_outputs_0_valid      (inputAll_3_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_3_ready                   ), //i
    .io_outputs_0_payload    (inputAll_3_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_3_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_3_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_3_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_4_fork (
    .io_input_valid          (inputAll_4_valid                      ), //i
    .io_input_ready          (inputAll_4_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_4_payload                    ), //i
    .io_outputs_0_valid      (inputAll_4_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_4_ready                   ), //i
    .io_outputs_0_payload    (inputAll_4_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_4_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_4_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_4_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_5_fork (
    .io_input_valid          (inputAll_5_valid                      ), //i
    .io_input_ready          (inputAll_5_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_5_payload                    ), //i
    .io_outputs_0_valid      (inputAll_5_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_5_ready                   ), //i
    .io_outputs_0_payload    (inputAll_5_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_5_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_5_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_5_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_6_fork (
    .io_input_valid          (inputAll_6_valid                      ), //i
    .io_input_ready          (inputAll_6_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_6_payload                    ), //i
    .io_outputs_0_valid      (inputAll_6_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_6_ready                   ), //i
    .io_outputs_0_payload    (inputAll_6_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_6_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_6_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_6_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_7_fork (
    .io_input_valid          (inputAll_7_valid                      ), //i
    .io_input_ready          (inputAll_7_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_7_payload                    ), //i
    .io_outputs_0_valid      (inputAll_7_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_7_ready                   ), //i
    .io_outputs_0_payload    (inputAll_7_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_7_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_7_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_7_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_8_fork (
    .io_input_valid          (inputAll_8_valid                      ), //i
    .io_input_ready          (inputAll_8_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_8_payload                    ), //i
    .io_outputs_0_valid      (inputAll_8_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_8_ready                   ), //i
    .io_outputs_0_payload    (inputAll_8_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_8_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_8_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_8_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_9_fork (
    .io_input_valid          (inputAll_9_valid                      ), //i
    .io_input_ready          (inputAll_9_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_9_payload                    ), //i
    .io_outputs_0_valid      (inputAll_9_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_9_ready                   ), //i
    .io_outputs_0_payload    (inputAll_9_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_9_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_9_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_9_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_10_fork (
    .io_input_valid          (inputAll_10_valid                      ), //i
    .io_input_ready          (inputAll_10_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_10_payload                    ), //i
    .io_outputs_0_valid      (inputAll_10_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_10_ready                   ), //i
    .io_outputs_0_payload    (inputAll_10_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_10_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_10_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_10_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_11_fork (
    .io_input_valid          (inputAll_11_valid                      ), //i
    .io_input_ready          (inputAll_11_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_11_payload                    ), //i
    .io_outputs_0_valid      (inputAll_11_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_11_ready                   ), //i
    .io_outputs_0_payload    (inputAll_11_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_11_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_11_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_11_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_12_fork (
    .io_input_valid          (inputAll_12_valid                      ), //i
    .io_input_ready          (inputAll_12_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_12_payload                    ), //i
    .io_outputs_0_valid      (inputAll_12_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_12_ready                   ), //i
    .io_outputs_0_payload    (inputAll_12_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_12_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_12_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_12_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_13_fork (
    .io_input_valid          (inputAll_13_valid                      ), //i
    .io_input_ready          (inputAll_13_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_13_payload                    ), //i
    .io_outputs_0_valid      (inputAll_13_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_13_ready                   ), //i
    .io_outputs_0_payload    (inputAll_13_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_13_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_13_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_13_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_14_fork (
    .io_input_valid          (inputAll_14_valid                      ), //i
    .io_input_ready          (inputAll_14_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_14_payload                    ), //i
    .io_outputs_0_valid      (inputAll_14_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_14_ready                   ), //i
    .io_outputs_0_payload    (inputAll_14_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_14_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_14_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_14_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_15_fork (
    .io_input_valid          (inputAll_15_valid                      ), //i
    .io_input_ready          (inputAll_15_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_15_payload                    ), //i
    .io_outputs_0_valid      (inputAll_15_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_15_ready                   ), //i
    .io_outputs_0_payload    (inputAll_15_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_15_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_15_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_15_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_16_fork (
    .io_input_valid          (inputAll_16_valid                      ), //i
    .io_input_ready          (inputAll_16_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_16_payload                    ), //i
    .io_outputs_0_valid      (inputAll_16_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_16_ready                   ), //i
    .io_outputs_0_payload    (inputAll_16_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_16_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_16_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_16_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_17_fork (
    .io_input_valid          (inputAll_17_valid                      ), //i
    .io_input_ready          (inputAll_17_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_17_payload                    ), //i
    .io_outputs_0_valid      (inputAll_17_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_17_ready                   ), //i
    .io_outputs_0_payload    (inputAll_17_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_17_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_17_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_17_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_18_fork (
    .io_input_valid          (inputAll_18_valid                      ), //i
    .io_input_ready          (inputAll_18_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_18_payload                    ), //i
    .io_outputs_0_valid      (inputAll_18_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_18_ready                   ), //i
    .io_outputs_0_payload    (inputAll_18_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_18_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_18_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_18_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_19_fork (
    .io_input_valid          (inputAll_19_valid                      ), //i
    .io_input_ready          (inputAll_19_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_19_payload                    ), //i
    .io_outputs_0_valid      (inputAll_19_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_19_ready                   ), //i
    .io_outputs_0_payload    (inputAll_19_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_19_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_19_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_19_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_20_fork (
    .io_input_valid          (inputAll_20_valid                      ), //i
    .io_input_ready          (inputAll_20_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_20_payload                    ), //i
    .io_outputs_0_valid      (inputAll_20_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_20_ready                   ), //i
    .io_outputs_0_payload    (inputAll_20_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_20_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_20_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_20_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_21_fork (
    .io_input_valid          (inputAll_21_valid                      ), //i
    .io_input_ready          (inputAll_21_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_21_payload                    ), //i
    .io_outputs_0_valid      (inputAll_21_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_21_ready                   ), //i
    .io_outputs_0_payload    (inputAll_21_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_21_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_21_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_21_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_22_fork (
    .io_input_valid          (inputAll_22_valid                      ), //i
    .io_input_ready          (inputAll_22_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_22_payload                    ), //i
    .io_outputs_0_valid      (inputAll_22_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_22_ready                   ), //i
    .io_outputs_0_payload    (inputAll_22_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_22_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_22_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_22_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_23_fork (
    .io_input_valid          (inputAll_23_valid                      ), //i
    .io_input_ready          (inputAll_23_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_23_payload                    ), //i
    .io_outputs_0_valid      (inputAll_23_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_23_ready                   ), //i
    .io_outputs_0_payload    (inputAll_23_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_23_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_23_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_23_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_24_fork (
    .io_input_valid          (inputAll_24_valid                      ), //i
    .io_input_ready          (inputAll_24_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_24_payload                    ), //i
    .io_outputs_0_valid      (inputAll_24_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_24_ready                   ), //i
    .io_outputs_0_payload    (inputAll_24_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_24_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_24_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_24_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_25_fork (
    .io_input_valid          (inputAll_25_valid                      ), //i
    .io_input_ready          (inputAll_25_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_25_payload                    ), //i
    .io_outputs_0_valid      (inputAll_25_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_25_ready                   ), //i
    .io_outputs_0_payload    (inputAll_25_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_25_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_25_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_25_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_26_fork (
    .io_input_valid          (inputAll_26_valid                      ), //i
    .io_input_ready          (inputAll_26_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_26_payload                    ), //i
    .io_outputs_0_valid      (inputAll_26_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_26_ready                   ), //i
    .io_outputs_0_payload    (inputAll_26_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_26_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_26_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_26_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_27_fork (
    .io_input_valid          (inputAll_27_valid                      ), //i
    .io_input_ready          (inputAll_27_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_27_payload                    ), //i
    .io_outputs_0_valid      (inputAll_27_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_27_ready                   ), //i
    .io_outputs_0_payload    (inputAll_27_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_27_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_27_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_27_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_28_fork (
    .io_input_valid          (inputAll_28_valid                      ), //i
    .io_input_ready          (inputAll_28_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_28_payload                    ), //i
    .io_outputs_0_valid      (inputAll_28_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_28_ready                   ), //i
    .io_outputs_0_payload    (inputAll_28_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_28_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_28_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_28_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_29_fork (
    .io_input_valid          (inputAll_29_valid                      ), //i
    .io_input_ready          (inputAll_29_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_29_payload                    ), //i
    .io_outputs_0_valid      (inputAll_29_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_29_ready                   ), //i
    .io_outputs_0_payload    (inputAll_29_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_29_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_29_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_29_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_30_fork (
    .io_input_valid          (inputAll_30_valid                      ), //i
    .io_input_ready          (inputAll_30_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_30_payload                    ), //i
    .io_outputs_0_valid      (inputAll_30_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_30_ready                   ), //i
    .io_outputs_0_payload    (inputAll_30_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_30_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_30_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_30_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_31_fork (
    .io_input_valid          (inputAll_31_valid                      ), //i
    .io_input_ready          (inputAll_31_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_31_payload                    ), //i
    .io_outputs_0_valid      (inputAll_31_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_31_ready                   ), //i
    .io_outputs_0_payload    (inputAll_31_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_31_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_31_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_31_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_32_fork (
    .io_input_valid          (inputAll_32_valid                      ), //i
    .io_input_ready          (inputAll_32_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_32_payload                    ), //i
    .io_outputs_0_valid      (inputAll_32_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_32_ready                   ), //i
    .io_outputs_0_payload    (inputAll_32_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_32_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_32_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_32_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_33_fork (
    .io_input_valid          (inputAll_33_valid                      ), //i
    .io_input_ready          (inputAll_33_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_33_payload                    ), //i
    .io_outputs_0_valid      (inputAll_33_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_33_ready                   ), //i
    .io_outputs_0_payload    (inputAll_33_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_33_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_33_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_33_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_34_fork (
    .io_input_valid          (inputAll_34_valid                      ), //i
    .io_input_ready          (inputAll_34_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_34_payload                    ), //i
    .io_outputs_0_valid      (inputAll_34_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_34_ready                   ), //i
    .io_outputs_0_payload    (inputAll_34_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_34_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_34_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_34_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_35_fork (
    .io_input_valid          (inputAll_35_valid                      ), //i
    .io_input_ready          (inputAll_35_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_35_payload                    ), //i
    .io_outputs_0_valid      (inputAll_35_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_35_ready                   ), //i
    .io_outputs_0_payload    (inputAll_35_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_35_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_35_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_35_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_36_fork (
    .io_input_valid          (inputAll_36_valid                      ), //i
    .io_input_ready          (inputAll_36_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_36_payload                    ), //i
    .io_outputs_0_valid      (inputAll_36_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_36_ready                   ), //i
    .io_outputs_0_payload    (inputAll_36_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_36_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_36_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_36_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_37_fork (
    .io_input_valid          (inputAll_37_valid                      ), //i
    .io_input_ready          (inputAll_37_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_37_payload                    ), //i
    .io_outputs_0_valid      (inputAll_37_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_37_ready                   ), //i
    .io_outputs_0_payload    (inputAll_37_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_37_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_37_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_37_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_38_fork (
    .io_input_valid          (inputAll_38_valid                      ), //i
    .io_input_ready          (inputAll_38_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_38_payload                    ), //i
    .io_outputs_0_valid      (inputAll_38_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_38_ready                   ), //i
    .io_outputs_0_payload    (inputAll_38_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_38_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_38_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_38_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_39_fork (
    .io_input_valid          (inputAll_39_valid                      ), //i
    .io_input_ready          (inputAll_39_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_39_payload                    ), //i
    .io_outputs_0_valid      (inputAll_39_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_39_ready                   ), //i
    .io_outputs_0_payload    (inputAll_39_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_39_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_39_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_39_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_40_fork (
    .io_input_valid          (inputAll_40_valid                      ), //i
    .io_input_ready          (inputAll_40_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_40_payload                    ), //i
    .io_outputs_0_valid      (inputAll_40_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_40_ready                   ), //i
    .io_outputs_0_payload    (inputAll_40_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_40_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_40_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_40_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_41_fork (
    .io_input_valid          (inputAll_41_valid                      ), //i
    .io_input_ready          (inputAll_41_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_41_payload                    ), //i
    .io_outputs_0_valid      (inputAll_41_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_41_ready                   ), //i
    .io_outputs_0_payload    (inputAll_41_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_41_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_41_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_41_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_42_fork (
    .io_input_valid          (inputAll_42_valid                      ), //i
    .io_input_ready          (inputAll_42_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_42_payload                    ), //i
    .io_outputs_0_valid      (inputAll_42_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_42_ready                   ), //i
    .io_outputs_0_payload    (inputAll_42_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_42_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_42_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_42_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_43_fork (
    .io_input_valid          (inputAll_43_valid                      ), //i
    .io_input_ready          (inputAll_43_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_43_payload                    ), //i
    .io_outputs_0_valid      (inputAll_43_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_43_ready                   ), //i
    .io_outputs_0_payload    (inputAll_43_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_43_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_43_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_43_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_44_fork (
    .io_input_valid          (inputAll_44_valid                      ), //i
    .io_input_ready          (inputAll_44_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_44_payload                    ), //i
    .io_outputs_0_valid      (inputAll_44_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_44_ready                   ), //i
    .io_outputs_0_payload    (inputAll_44_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_44_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_44_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_44_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_45_fork (
    .io_input_valid          (inputAll_45_valid                      ), //i
    .io_input_ready          (inputAll_45_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_45_payload                    ), //i
    .io_outputs_0_valid      (inputAll_45_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_45_ready                   ), //i
    .io_outputs_0_payload    (inputAll_45_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_45_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_45_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_45_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_46_fork (
    .io_input_valid          (inputAll_46_valid                      ), //i
    .io_input_ready          (inputAll_46_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_46_payload                    ), //i
    .io_outputs_0_valid      (inputAll_46_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_46_ready                   ), //i
    .io_outputs_0_payload    (inputAll_46_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_46_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_46_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_46_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_47_fork (
    .io_input_valid          (inputAll_47_valid                      ), //i
    .io_input_ready          (inputAll_47_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_47_payload                    ), //i
    .io_outputs_0_valid      (inputAll_47_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_47_ready                   ), //i
    .io_outputs_0_payload    (inputAll_47_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_47_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_47_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_47_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_48_fork (
    .io_input_valid          (inputAll_48_valid                      ), //i
    .io_input_ready          (inputAll_48_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_48_payload                    ), //i
    .io_outputs_0_valid      (inputAll_48_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_48_ready                   ), //i
    .io_outputs_0_payload    (inputAll_48_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_48_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_48_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_48_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_49_fork (
    .io_input_valid          (inputAll_49_valid                      ), //i
    .io_input_ready          (inputAll_49_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_49_payload                    ), //i
    .io_outputs_0_valid      (inputAll_49_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_49_ready                   ), //i
    .io_outputs_0_payload    (inputAll_49_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_49_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_49_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_49_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_50_fork (
    .io_input_valid          (inputAll_50_valid                      ), //i
    .io_input_ready          (inputAll_50_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_50_payload                    ), //i
    .io_outputs_0_valid      (inputAll_50_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_50_ready                   ), //i
    .io_outputs_0_payload    (inputAll_50_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_50_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_50_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_50_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_51_fork (
    .io_input_valid          (inputAll_51_valid                      ), //i
    .io_input_ready          (inputAll_51_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_51_payload                    ), //i
    .io_outputs_0_valid      (inputAll_51_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_51_ready                   ), //i
    .io_outputs_0_payload    (inputAll_51_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_51_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_51_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_51_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_52_fork (
    .io_input_valid          (inputAll_52_valid                      ), //i
    .io_input_ready          (inputAll_52_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_52_payload                    ), //i
    .io_outputs_0_valid      (inputAll_52_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_52_ready                   ), //i
    .io_outputs_0_payload    (inputAll_52_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_52_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_52_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_52_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_53_fork (
    .io_input_valid          (inputAll_53_valid                      ), //i
    .io_input_ready          (inputAll_53_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_53_payload                    ), //i
    .io_outputs_0_valid      (inputAll_53_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_53_ready                   ), //i
    .io_outputs_0_payload    (inputAll_53_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_53_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_53_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_53_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_54_fork (
    .io_input_valid          (inputAll_54_valid                      ), //i
    .io_input_ready          (inputAll_54_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_54_payload                    ), //i
    .io_outputs_0_valid      (inputAll_54_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_54_ready                   ), //i
    .io_outputs_0_payload    (inputAll_54_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_54_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_54_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_54_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_55_fork (
    .io_input_valid          (inputAll_55_valid                      ), //i
    .io_input_ready          (inputAll_55_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_55_payload                    ), //i
    .io_outputs_0_valid      (inputAll_55_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_55_ready                   ), //i
    .io_outputs_0_payload    (inputAll_55_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_55_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_55_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_55_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_56_fork (
    .io_input_valid          (inputAll_56_valid                      ), //i
    .io_input_ready          (inputAll_56_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_56_payload                    ), //i
    .io_outputs_0_valid      (inputAll_56_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_56_ready                   ), //i
    .io_outputs_0_payload    (inputAll_56_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_56_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_56_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_56_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_57_fork (
    .io_input_valid          (inputAll_57_valid                      ), //i
    .io_input_ready          (inputAll_57_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_57_payload                    ), //i
    .io_outputs_0_valid      (inputAll_57_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_57_ready                   ), //i
    .io_outputs_0_payload    (inputAll_57_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_57_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_57_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_57_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_58_fork (
    .io_input_valid          (inputAll_58_valid                      ), //i
    .io_input_ready          (inputAll_58_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_58_payload                    ), //i
    .io_outputs_0_valid      (inputAll_58_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_58_ready                   ), //i
    .io_outputs_0_payload    (inputAll_58_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_58_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_58_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_58_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_59_fork (
    .io_input_valid          (inputAll_59_valid                      ), //i
    .io_input_ready          (inputAll_59_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_59_payload                    ), //i
    .io_outputs_0_valid      (inputAll_59_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_59_ready                   ), //i
    .io_outputs_0_payload    (inputAll_59_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_59_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_59_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_59_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_60_fork (
    .io_input_valid          (inputAll_60_valid                      ), //i
    .io_input_ready          (inputAll_60_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_60_payload                    ), //i
    .io_outputs_0_valid      (inputAll_60_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_60_ready                   ), //i
    .io_outputs_0_payload    (inputAll_60_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_60_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_60_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_60_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_61_fork (
    .io_input_valid          (inputAll_61_valid                      ), //i
    .io_input_ready          (inputAll_61_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_61_payload                    ), //i
    .io_outputs_0_valid      (inputAll_61_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_61_ready                   ), //i
    .io_outputs_0_payload    (inputAll_61_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_61_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_61_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_61_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_62_fork (
    .io_input_valid          (inputAll_62_valid                      ), //i
    .io_input_ready          (inputAll_62_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_62_payload                    ), //i
    .io_outputs_0_valid      (inputAll_62_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_62_ready                   ), //i
    .io_outputs_0_payload    (inputAll_62_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_62_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_62_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_62_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_63_fork (
    .io_input_valid          (inputAll_63_valid                      ), //i
    .io_input_ready          (inputAll_63_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_63_payload                    ), //i
    .io_outputs_0_valid      (inputAll_63_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_63_ready                   ), //i
    .io_outputs_0_payload    (inputAll_63_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_63_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_63_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_63_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_64_fork (
    .io_input_valid          (inputAll_64_valid                      ), //i
    .io_input_ready          (inputAll_64_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_64_payload                    ), //i
    .io_outputs_0_valid      (inputAll_64_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_63_ready                   ), //i
    .io_outputs_0_payload    (inputAll_64_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_64_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_64_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_64_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_65_fork (
    .io_input_valid          (inputAll_65_valid                      ), //i
    .io_input_ready          (inputAll_65_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_65_payload                    ), //i
    .io_outputs_0_valid      (inputAll_65_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_62_ready                   ), //i
    .io_outputs_0_payload    (inputAll_65_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_65_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_65_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_65_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_66_fork (
    .io_input_valid          (inputAll_66_valid                      ), //i
    .io_input_ready          (inputAll_66_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_66_payload                    ), //i
    .io_outputs_0_valid      (inputAll_66_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_61_ready                   ), //i
    .io_outputs_0_payload    (inputAll_66_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_66_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_66_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_66_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_67_fork (
    .io_input_valid          (inputAll_67_valid                      ), //i
    .io_input_ready          (inputAll_67_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_67_payload                    ), //i
    .io_outputs_0_valid      (inputAll_67_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_60_ready                   ), //i
    .io_outputs_0_payload    (inputAll_67_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_67_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_67_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_67_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_68_fork (
    .io_input_valid          (inputAll_68_valid                      ), //i
    .io_input_ready          (inputAll_68_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_68_payload                    ), //i
    .io_outputs_0_valid      (inputAll_68_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_59_ready                   ), //i
    .io_outputs_0_payload    (inputAll_68_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_68_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_68_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_68_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_69_fork (
    .io_input_valid          (inputAll_69_valid                      ), //i
    .io_input_ready          (inputAll_69_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_69_payload                    ), //i
    .io_outputs_0_valid      (inputAll_69_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_58_ready                   ), //i
    .io_outputs_0_payload    (inputAll_69_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_69_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_69_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_69_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_70_fork (
    .io_input_valid          (inputAll_70_valid                      ), //i
    .io_input_ready          (inputAll_70_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_70_payload                    ), //i
    .io_outputs_0_valid      (inputAll_70_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_57_ready                   ), //i
    .io_outputs_0_payload    (inputAll_70_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_70_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_70_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_70_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_71_fork (
    .io_input_valid          (inputAll_71_valid                      ), //i
    .io_input_ready          (inputAll_71_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_71_payload                    ), //i
    .io_outputs_0_valid      (inputAll_71_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_56_ready                   ), //i
    .io_outputs_0_payload    (inputAll_71_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_71_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_71_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_71_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_72_fork (
    .io_input_valid          (inputAll_72_valid                      ), //i
    .io_input_ready          (inputAll_72_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_72_payload                    ), //i
    .io_outputs_0_valid      (inputAll_72_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_55_ready                   ), //i
    .io_outputs_0_payload    (inputAll_72_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_72_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_72_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_72_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_73_fork (
    .io_input_valid          (inputAll_73_valid                      ), //i
    .io_input_ready          (inputAll_73_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_73_payload                    ), //i
    .io_outputs_0_valid      (inputAll_73_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_54_ready                   ), //i
    .io_outputs_0_payload    (inputAll_73_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_73_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_73_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_73_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_74_fork (
    .io_input_valid          (inputAll_74_valid                      ), //i
    .io_input_ready          (inputAll_74_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_74_payload                    ), //i
    .io_outputs_0_valid      (inputAll_74_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_53_ready                   ), //i
    .io_outputs_0_payload    (inputAll_74_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_74_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_74_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_74_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_75_fork (
    .io_input_valid          (inputAll_75_valid                      ), //i
    .io_input_ready          (inputAll_75_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_75_payload                    ), //i
    .io_outputs_0_valid      (inputAll_75_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_52_ready                   ), //i
    .io_outputs_0_payload    (inputAll_75_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_75_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_75_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_75_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_76_fork (
    .io_input_valid          (inputAll_76_valid                      ), //i
    .io_input_ready          (inputAll_76_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_76_payload                    ), //i
    .io_outputs_0_valid      (inputAll_76_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_51_ready                   ), //i
    .io_outputs_0_payload    (inputAll_76_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_76_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_76_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_76_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_77_fork (
    .io_input_valid          (inputAll_77_valid                      ), //i
    .io_input_ready          (inputAll_77_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_77_payload                    ), //i
    .io_outputs_0_valid      (inputAll_77_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_50_ready                   ), //i
    .io_outputs_0_payload    (inputAll_77_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_77_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_77_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_77_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_78_fork (
    .io_input_valid          (inputAll_78_valid                      ), //i
    .io_input_ready          (inputAll_78_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_78_payload                    ), //i
    .io_outputs_0_valid      (inputAll_78_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_49_ready                   ), //i
    .io_outputs_0_payload    (inputAll_78_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_78_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_78_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_78_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_79_fork (
    .io_input_valid          (inputAll_79_valid                      ), //i
    .io_input_ready          (inputAll_79_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_79_payload                    ), //i
    .io_outputs_0_valid      (inputAll_79_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_48_ready                   ), //i
    .io_outputs_0_payload    (inputAll_79_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_79_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_79_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_79_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_80_fork (
    .io_input_valid          (inputAll_80_valid                      ), //i
    .io_input_ready          (inputAll_80_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_80_payload                    ), //i
    .io_outputs_0_valid      (inputAll_80_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_47_ready                   ), //i
    .io_outputs_0_payload    (inputAll_80_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_80_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_80_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_80_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_81_fork (
    .io_input_valid          (inputAll_81_valid                      ), //i
    .io_input_ready          (inputAll_81_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_81_payload                    ), //i
    .io_outputs_0_valid      (inputAll_81_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_46_ready                   ), //i
    .io_outputs_0_payload    (inputAll_81_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_81_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_81_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_81_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_82_fork (
    .io_input_valid          (inputAll_82_valid                      ), //i
    .io_input_ready          (inputAll_82_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_82_payload                    ), //i
    .io_outputs_0_valid      (inputAll_82_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_45_ready                   ), //i
    .io_outputs_0_payload    (inputAll_82_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_82_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_82_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_82_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_83_fork (
    .io_input_valid          (inputAll_83_valid                      ), //i
    .io_input_ready          (inputAll_83_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_83_payload                    ), //i
    .io_outputs_0_valid      (inputAll_83_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_44_ready                   ), //i
    .io_outputs_0_payload    (inputAll_83_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_83_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_83_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_83_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_84_fork (
    .io_input_valid          (inputAll_84_valid                      ), //i
    .io_input_ready          (inputAll_84_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_84_payload                    ), //i
    .io_outputs_0_valid      (inputAll_84_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_43_ready                   ), //i
    .io_outputs_0_payload    (inputAll_84_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_84_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_84_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_84_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_85_fork (
    .io_input_valid          (inputAll_85_valid                      ), //i
    .io_input_ready          (inputAll_85_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_85_payload                    ), //i
    .io_outputs_0_valid      (inputAll_85_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_42_ready                   ), //i
    .io_outputs_0_payload    (inputAll_85_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_85_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_85_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_85_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_86_fork (
    .io_input_valid          (inputAll_86_valid                      ), //i
    .io_input_ready          (inputAll_86_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_86_payload                    ), //i
    .io_outputs_0_valid      (inputAll_86_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_41_ready                   ), //i
    .io_outputs_0_payload    (inputAll_86_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_86_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_86_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_86_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_87_fork (
    .io_input_valid          (inputAll_87_valid                      ), //i
    .io_input_ready          (inputAll_87_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_87_payload                    ), //i
    .io_outputs_0_valid      (inputAll_87_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_40_ready                   ), //i
    .io_outputs_0_payload    (inputAll_87_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_87_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_87_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_87_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_88_fork (
    .io_input_valid          (inputAll_88_valid                      ), //i
    .io_input_ready          (inputAll_88_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_88_payload                    ), //i
    .io_outputs_0_valid      (inputAll_88_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_39_ready                   ), //i
    .io_outputs_0_payload    (inputAll_88_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_88_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_88_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_88_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_89_fork (
    .io_input_valid          (inputAll_89_valid                      ), //i
    .io_input_ready          (inputAll_89_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_89_payload                    ), //i
    .io_outputs_0_valid      (inputAll_89_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_38_ready                   ), //i
    .io_outputs_0_payload    (inputAll_89_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_89_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_89_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_89_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_90_fork (
    .io_input_valid          (inputAll_90_valid                      ), //i
    .io_input_ready          (inputAll_90_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_90_payload                    ), //i
    .io_outputs_0_valid      (inputAll_90_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_37_ready                   ), //i
    .io_outputs_0_payload    (inputAll_90_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_90_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_90_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_90_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_91_fork (
    .io_input_valid          (inputAll_91_valid                      ), //i
    .io_input_ready          (inputAll_91_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_91_payload                    ), //i
    .io_outputs_0_valid      (inputAll_91_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_36_ready                   ), //i
    .io_outputs_0_payload    (inputAll_91_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_91_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_91_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_91_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_92_fork (
    .io_input_valid          (inputAll_92_valid                      ), //i
    .io_input_ready          (inputAll_92_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_92_payload                    ), //i
    .io_outputs_0_valid      (inputAll_92_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_35_ready                   ), //i
    .io_outputs_0_payload    (inputAll_92_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_92_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_92_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_92_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_93_fork (
    .io_input_valid          (inputAll_93_valid                      ), //i
    .io_input_ready          (inputAll_93_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_93_payload                    ), //i
    .io_outputs_0_valid      (inputAll_93_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_34_ready                   ), //i
    .io_outputs_0_payload    (inputAll_93_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_93_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_93_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_93_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_94_fork (
    .io_input_valid          (inputAll_94_valid                      ), //i
    .io_input_ready          (inputAll_94_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_94_payload                    ), //i
    .io_outputs_0_valid      (inputAll_94_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_33_ready                   ), //i
    .io_outputs_0_payload    (inputAll_94_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_94_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_94_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_94_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_95_fork (
    .io_input_valid          (inputAll_95_valid                      ), //i
    .io_input_ready          (inputAll_95_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_95_payload                    ), //i
    .io_outputs_0_valid      (inputAll_95_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_32_ready                   ), //i
    .io_outputs_0_payload    (inputAll_95_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_95_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_95_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_95_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_96_fork (
    .io_input_valid          (inputAll_96_valid                      ), //i
    .io_input_ready          (inputAll_96_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_96_payload                    ), //i
    .io_outputs_0_valid      (inputAll_96_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_31_ready                   ), //i
    .io_outputs_0_payload    (inputAll_96_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_96_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_96_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_96_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_97_fork (
    .io_input_valid          (inputAll_97_valid                      ), //i
    .io_input_ready          (inputAll_97_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_97_payload                    ), //i
    .io_outputs_0_valid      (inputAll_97_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_30_ready                   ), //i
    .io_outputs_0_payload    (inputAll_97_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_97_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_97_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_97_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_98_fork (
    .io_input_valid          (inputAll_98_valid                      ), //i
    .io_input_ready          (inputAll_98_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_98_payload                    ), //i
    .io_outputs_0_valid      (inputAll_98_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_29_ready                   ), //i
    .io_outputs_0_payload    (inputAll_98_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_98_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_98_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_98_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_99_fork (
    .io_input_valid          (inputAll_99_valid                      ), //i
    .io_input_ready          (inputAll_99_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_99_payload                    ), //i
    .io_outputs_0_valid      (inputAll_99_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_28_ready                   ), //i
    .io_outputs_0_payload    (inputAll_99_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_99_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_99_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_99_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_100_fork (
    .io_input_valid          (inputAll_100_valid                      ), //i
    .io_input_ready          (inputAll_100_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_100_payload                    ), //i
    .io_outputs_0_valid      (inputAll_100_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_27_ready                    ), //i
    .io_outputs_0_payload    (inputAll_100_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_100_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_100_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_100_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_101_fork (
    .io_input_valid          (inputAll_101_valid                      ), //i
    .io_input_ready          (inputAll_101_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_101_payload                    ), //i
    .io_outputs_0_valid      (inputAll_101_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_26_ready                    ), //i
    .io_outputs_0_payload    (inputAll_101_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_101_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_101_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_101_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_102_fork (
    .io_input_valid          (inputAll_102_valid                      ), //i
    .io_input_ready          (inputAll_102_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_102_payload                    ), //i
    .io_outputs_0_valid      (inputAll_102_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_25_ready                    ), //i
    .io_outputs_0_payload    (inputAll_102_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_102_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_102_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_102_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_103_fork (
    .io_input_valid          (inputAll_103_valid                      ), //i
    .io_input_ready          (inputAll_103_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_103_payload                    ), //i
    .io_outputs_0_valid      (inputAll_103_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_24_ready                    ), //i
    .io_outputs_0_payload    (inputAll_103_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_103_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_103_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_103_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_104_fork (
    .io_input_valid          (inputAll_104_valid                      ), //i
    .io_input_ready          (inputAll_104_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_104_payload                    ), //i
    .io_outputs_0_valid      (inputAll_104_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_23_ready                    ), //i
    .io_outputs_0_payload    (inputAll_104_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_104_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_104_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_104_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_105_fork (
    .io_input_valid          (inputAll_105_valid                      ), //i
    .io_input_ready          (inputAll_105_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_105_payload                    ), //i
    .io_outputs_0_valid      (inputAll_105_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_22_ready                    ), //i
    .io_outputs_0_payload    (inputAll_105_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_105_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_105_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_105_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_106_fork (
    .io_input_valid          (inputAll_106_valid                      ), //i
    .io_input_ready          (inputAll_106_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_106_payload                    ), //i
    .io_outputs_0_valid      (inputAll_106_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_21_ready                    ), //i
    .io_outputs_0_payload    (inputAll_106_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_106_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_106_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_106_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_107_fork (
    .io_input_valid          (inputAll_107_valid                      ), //i
    .io_input_ready          (inputAll_107_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_107_payload                    ), //i
    .io_outputs_0_valid      (inputAll_107_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_20_ready                    ), //i
    .io_outputs_0_payload    (inputAll_107_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_107_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_107_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_107_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_108_fork (
    .io_input_valid          (inputAll_108_valid                      ), //i
    .io_input_ready          (inputAll_108_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_108_payload                    ), //i
    .io_outputs_0_valid      (inputAll_108_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_19_ready                    ), //i
    .io_outputs_0_payload    (inputAll_108_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_108_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_108_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_108_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_109_fork (
    .io_input_valid          (inputAll_109_valid                      ), //i
    .io_input_ready          (inputAll_109_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_109_payload                    ), //i
    .io_outputs_0_valid      (inputAll_109_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_18_ready                    ), //i
    .io_outputs_0_payload    (inputAll_109_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_109_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_109_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_109_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_110_fork (
    .io_input_valid          (inputAll_110_valid                      ), //i
    .io_input_ready          (inputAll_110_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_110_payload                    ), //i
    .io_outputs_0_valid      (inputAll_110_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_17_ready                    ), //i
    .io_outputs_0_payload    (inputAll_110_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_110_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_110_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_110_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_111_fork (
    .io_input_valid          (inputAll_111_valid                      ), //i
    .io_input_ready          (inputAll_111_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_111_payload                    ), //i
    .io_outputs_0_valid      (inputAll_111_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_16_ready                    ), //i
    .io_outputs_0_payload    (inputAll_111_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_111_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_111_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_111_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_112_fork (
    .io_input_valid          (inputAll_112_valid                      ), //i
    .io_input_ready          (inputAll_112_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_112_payload                    ), //i
    .io_outputs_0_valid      (inputAll_112_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_15_ready                    ), //i
    .io_outputs_0_payload    (inputAll_112_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_112_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_112_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_112_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_113_fork (
    .io_input_valid          (inputAll_113_valid                      ), //i
    .io_input_ready          (inputAll_113_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_113_payload                    ), //i
    .io_outputs_0_valid      (inputAll_113_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_14_ready                    ), //i
    .io_outputs_0_payload    (inputAll_113_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_113_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_113_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_113_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_114_fork (
    .io_input_valid          (inputAll_114_valid                      ), //i
    .io_input_ready          (inputAll_114_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_114_payload                    ), //i
    .io_outputs_0_valid      (inputAll_114_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_13_ready                    ), //i
    .io_outputs_0_payload    (inputAll_114_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_114_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_114_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_114_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_115_fork (
    .io_input_valid          (inputAll_115_valid                      ), //i
    .io_input_ready          (inputAll_115_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_115_payload                    ), //i
    .io_outputs_0_valid      (inputAll_115_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_12_ready                    ), //i
    .io_outputs_0_payload    (inputAll_115_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_115_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_115_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_115_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_116_fork (
    .io_input_valid          (inputAll_116_valid                      ), //i
    .io_input_ready          (inputAll_116_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_116_payload                    ), //i
    .io_outputs_0_valid      (inputAll_116_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_11_ready                    ), //i
    .io_outputs_0_payload    (inputAll_116_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_116_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_116_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_116_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_117_fork (
    .io_input_valid          (inputAll_117_valid                      ), //i
    .io_input_ready          (inputAll_117_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_117_payload                    ), //i
    .io_outputs_0_valid      (inputAll_117_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_10_ready                    ), //i
    .io_outputs_0_payload    (inputAll_117_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_117_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_117_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_117_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_118_fork (
    .io_input_valid          (inputAll_118_valid                      ), //i
    .io_input_ready          (inputAll_118_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_118_payload                    ), //i
    .io_outputs_0_valid      (inputAll_118_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_9_ready                     ), //i
    .io_outputs_0_payload    (inputAll_118_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_118_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_118_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_118_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_119_fork (
    .io_input_valid          (inputAll_119_valid                      ), //i
    .io_input_ready          (inputAll_119_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_119_payload                    ), //i
    .io_outputs_0_valid      (inputAll_119_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_8_ready                     ), //i
    .io_outputs_0_payload    (inputAll_119_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_119_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_119_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_119_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_120_fork (
    .io_input_valid          (inputAll_120_valid                      ), //i
    .io_input_ready          (inputAll_120_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_120_payload                    ), //i
    .io_outputs_0_valid      (inputAll_120_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_7_ready                     ), //i
    .io_outputs_0_payload    (inputAll_120_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_120_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_120_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_120_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_121_fork (
    .io_input_valid          (inputAll_121_valid                      ), //i
    .io_input_ready          (inputAll_121_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_121_payload                    ), //i
    .io_outputs_0_valid      (inputAll_121_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_6_ready                     ), //i
    .io_outputs_0_payload    (inputAll_121_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_121_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_121_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_121_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_122_fork (
    .io_input_valid          (inputAll_122_valid                      ), //i
    .io_input_ready          (inputAll_122_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_122_payload                    ), //i
    .io_outputs_0_valid      (inputAll_122_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_5_ready                     ), //i
    .io_outputs_0_payload    (inputAll_122_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_122_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_122_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_122_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_123_fork (
    .io_input_valid          (inputAll_123_valid                      ), //i
    .io_input_ready          (inputAll_123_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_123_payload                    ), //i
    .io_outputs_0_valid      (inputAll_123_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_4_ready                     ), //i
    .io_outputs_0_payload    (inputAll_123_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_123_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_123_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_123_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_124_fork (
    .io_input_valid          (inputAll_124_valid                      ), //i
    .io_input_ready          (inputAll_124_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_124_payload                    ), //i
    .io_outputs_0_valid      (inputAll_124_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_3_ready                     ), //i
    .io_outputs_0_payload    (inputAll_124_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_124_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_124_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_124_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_125_fork (
    .io_input_valid          (inputAll_125_valid                      ), //i
    .io_input_ready          (inputAll_125_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_125_payload                    ), //i
    .io_outputs_0_valid      (inputAll_125_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_2_ready                     ), //i
    .io_outputs_0_payload    (inputAll_125_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_125_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_125_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_125_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_126_fork (
    .io_input_valid          (inputAll_126_valid                      ), //i
    .io_input_ready          (inputAll_126_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_126_payload                    ), //i
    .io_outputs_0_valid      (inputAll_126_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_1_ready                     ), //i
    .io_outputs_0_payload    (inputAll_126_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_126_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_126_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_126_fork_io_outputs_1_payload  )  //o
  );
  StreamFork inputAll_127_fork (
    .io_input_valid          (inputAll_127_valid                      ), //i
    .io_input_ready          (inputAll_127_fork_io_input_ready        ), //o
    .io_input_payload        (inputAll_127_payload                    ), //i
    .io_outputs_0_valid      (inputAll_127_fork_io_outputs_0_valid    ), //o
    .io_outputs_0_ready      (mulResGroup_0_ready                     ), //i
    .io_outputs_0_payload    (inputAll_127_fork_io_outputs_0_payload  ), //o
    .io_outputs_1_valid      (inputAll_127_fork_io_outputs_1_valid    ), //o
    .io_outputs_1_ready      (inputAll_127_fork_io_outputs_1_ready    ), //i
    .io_outputs_1_payload    (inputAll_127_fork_io_outputs_1_payload  )  //o
  );
  assign inputAll_0_ready = inputAll_0_fork_io_input_ready;
  always @(*) begin
    inputAll_0_fork_io_outputs_1_ready = inputAll_0_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342) begin
      inputAll_0_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! inputAll_0_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_0_fork_io_outputs_1_m2sPipe_valid = inputAll_0_fork_io_outputs_1_rValid;
  assign inputAll_0_fork_io_outputs_1_m2sPipe_payload = inputAll_0_fork_io_outputs_1_rData;
  assign inputAll_1_ready = inputAll_1_fork_io_input_ready;
  always @(*) begin
    inputAll_1_fork_io_outputs_1_ready = inputAll_1_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      inputAll_1_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! inputAll_1_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_1_fork_io_outputs_1_m2sPipe_valid = inputAll_1_fork_io_outputs_1_rValid;
  assign inputAll_1_fork_io_outputs_1_m2sPipe_payload = inputAll_1_fork_io_outputs_1_rData;
  assign inputAll_2_ready = inputAll_2_fork_io_input_ready;
  always @(*) begin
    inputAll_2_fork_io_outputs_1_ready = inputAll_2_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      inputAll_2_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! inputAll_2_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_2_fork_io_outputs_1_m2sPipe_valid = inputAll_2_fork_io_outputs_1_rValid;
  assign inputAll_2_fork_io_outputs_1_m2sPipe_payload = inputAll_2_fork_io_outputs_1_rData;
  assign inputAll_3_ready = inputAll_3_fork_io_input_ready;
  always @(*) begin
    inputAll_3_fork_io_outputs_1_ready = inputAll_3_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_3) begin
      inputAll_3_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! inputAll_3_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_3_fork_io_outputs_1_m2sPipe_valid = inputAll_3_fork_io_outputs_1_rValid;
  assign inputAll_3_fork_io_outputs_1_m2sPipe_payload = inputAll_3_fork_io_outputs_1_rData;
  assign inputAll_4_ready = inputAll_4_fork_io_input_ready;
  always @(*) begin
    inputAll_4_fork_io_outputs_1_ready = inputAll_4_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_4) begin
      inputAll_4_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! inputAll_4_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_4_fork_io_outputs_1_m2sPipe_valid = inputAll_4_fork_io_outputs_1_rValid;
  assign inputAll_4_fork_io_outputs_1_m2sPipe_payload = inputAll_4_fork_io_outputs_1_rData;
  assign inputAll_5_ready = inputAll_5_fork_io_input_ready;
  always @(*) begin
    inputAll_5_fork_io_outputs_1_ready = inputAll_5_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_5) begin
      inputAll_5_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! inputAll_5_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_5_fork_io_outputs_1_m2sPipe_valid = inputAll_5_fork_io_outputs_1_rValid;
  assign inputAll_5_fork_io_outputs_1_m2sPipe_payload = inputAll_5_fork_io_outputs_1_rData;
  assign inputAll_6_ready = inputAll_6_fork_io_input_ready;
  always @(*) begin
    inputAll_6_fork_io_outputs_1_ready = inputAll_6_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_6) begin
      inputAll_6_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_6 = (! inputAll_6_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_6_fork_io_outputs_1_m2sPipe_valid = inputAll_6_fork_io_outputs_1_rValid;
  assign inputAll_6_fork_io_outputs_1_m2sPipe_payload = inputAll_6_fork_io_outputs_1_rData;
  assign inputAll_7_ready = inputAll_7_fork_io_input_ready;
  always @(*) begin
    inputAll_7_fork_io_outputs_1_ready = inputAll_7_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_7) begin
      inputAll_7_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_7 = (! inputAll_7_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_7_fork_io_outputs_1_m2sPipe_valid = inputAll_7_fork_io_outputs_1_rValid;
  assign inputAll_7_fork_io_outputs_1_m2sPipe_payload = inputAll_7_fork_io_outputs_1_rData;
  assign inputAll_8_ready = inputAll_8_fork_io_input_ready;
  always @(*) begin
    inputAll_8_fork_io_outputs_1_ready = inputAll_8_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_8) begin
      inputAll_8_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_8 = (! inputAll_8_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_8_fork_io_outputs_1_m2sPipe_valid = inputAll_8_fork_io_outputs_1_rValid;
  assign inputAll_8_fork_io_outputs_1_m2sPipe_payload = inputAll_8_fork_io_outputs_1_rData;
  assign inputAll_9_ready = inputAll_9_fork_io_input_ready;
  always @(*) begin
    inputAll_9_fork_io_outputs_1_ready = inputAll_9_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_9) begin
      inputAll_9_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_9 = (! inputAll_9_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_9_fork_io_outputs_1_m2sPipe_valid = inputAll_9_fork_io_outputs_1_rValid;
  assign inputAll_9_fork_io_outputs_1_m2sPipe_payload = inputAll_9_fork_io_outputs_1_rData;
  assign inputAll_10_ready = inputAll_10_fork_io_input_ready;
  always @(*) begin
    inputAll_10_fork_io_outputs_1_ready = inputAll_10_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_10) begin
      inputAll_10_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_10 = (! inputAll_10_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_10_fork_io_outputs_1_m2sPipe_valid = inputAll_10_fork_io_outputs_1_rValid;
  assign inputAll_10_fork_io_outputs_1_m2sPipe_payload = inputAll_10_fork_io_outputs_1_rData;
  assign inputAll_11_ready = inputAll_11_fork_io_input_ready;
  always @(*) begin
    inputAll_11_fork_io_outputs_1_ready = inputAll_11_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_11) begin
      inputAll_11_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_11 = (! inputAll_11_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_11_fork_io_outputs_1_m2sPipe_valid = inputAll_11_fork_io_outputs_1_rValid;
  assign inputAll_11_fork_io_outputs_1_m2sPipe_payload = inputAll_11_fork_io_outputs_1_rData;
  assign inputAll_12_ready = inputAll_12_fork_io_input_ready;
  always @(*) begin
    inputAll_12_fork_io_outputs_1_ready = inputAll_12_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_12) begin
      inputAll_12_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_12 = (! inputAll_12_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_12_fork_io_outputs_1_m2sPipe_valid = inputAll_12_fork_io_outputs_1_rValid;
  assign inputAll_12_fork_io_outputs_1_m2sPipe_payload = inputAll_12_fork_io_outputs_1_rData;
  assign inputAll_13_ready = inputAll_13_fork_io_input_ready;
  always @(*) begin
    inputAll_13_fork_io_outputs_1_ready = inputAll_13_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_13) begin
      inputAll_13_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_13 = (! inputAll_13_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_13_fork_io_outputs_1_m2sPipe_valid = inputAll_13_fork_io_outputs_1_rValid;
  assign inputAll_13_fork_io_outputs_1_m2sPipe_payload = inputAll_13_fork_io_outputs_1_rData;
  assign inputAll_14_ready = inputAll_14_fork_io_input_ready;
  always @(*) begin
    inputAll_14_fork_io_outputs_1_ready = inputAll_14_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_14) begin
      inputAll_14_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_14 = (! inputAll_14_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_14_fork_io_outputs_1_m2sPipe_valid = inputAll_14_fork_io_outputs_1_rValid;
  assign inputAll_14_fork_io_outputs_1_m2sPipe_payload = inputAll_14_fork_io_outputs_1_rData;
  assign inputAll_15_ready = inputAll_15_fork_io_input_ready;
  always @(*) begin
    inputAll_15_fork_io_outputs_1_ready = inputAll_15_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_15) begin
      inputAll_15_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_15 = (! inputAll_15_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_15_fork_io_outputs_1_m2sPipe_valid = inputAll_15_fork_io_outputs_1_rValid;
  assign inputAll_15_fork_io_outputs_1_m2sPipe_payload = inputAll_15_fork_io_outputs_1_rData;
  assign inputAll_16_ready = inputAll_16_fork_io_input_ready;
  always @(*) begin
    inputAll_16_fork_io_outputs_1_ready = inputAll_16_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_16) begin
      inputAll_16_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_16 = (! inputAll_16_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_16_fork_io_outputs_1_m2sPipe_valid = inputAll_16_fork_io_outputs_1_rValid;
  assign inputAll_16_fork_io_outputs_1_m2sPipe_payload = inputAll_16_fork_io_outputs_1_rData;
  assign inputAll_17_ready = inputAll_17_fork_io_input_ready;
  always @(*) begin
    inputAll_17_fork_io_outputs_1_ready = inputAll_17_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_17) begin
      inputAll_17_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_17 = (! inputAll_17_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_17_fork_io_outputs_1_m2sPipe_valid = inputAll_17_fork_io_outputs_1_rValid;
  assign inputAll_17_fork_io_outputs_1_m2sPipe_payload = inputAll_17_fork_io_outputs_1_rData;
  assign inputAll_18_ready = inputAll_18_fork_io_input_ready;
  always @(*) begin
    inputAll_18_fork_io_outputs_1_ready = inputAll_18_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_18) begin
      inputAll_18_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_18 = (! inputAll_18_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_18_fork_io_outputs_1_m2sPipe_valid = inputAll_18_fork_io_outputs_1_rValid;
  assign inputAll_18_fork_io_outputs_1_m2sPipe_payload = inputAll_18_fork_io_outputs_1_rData;
  assign inputAll_19_ready = inputAll_19_fork_io_input_ready;
  always @(*) begin
    inputAll_19_fork_io_outputs_1_ready = inputAll_19_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_19) begin
      inputAll_19_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_19 = (! inputAll_19_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_19_fork_io_outputs_1_m2sPipe_valid = inputAll_19_fork_io_outputs_1_rValid;
  assign inputAll_19_fork_io_outputs_1_m2sPipe_payload = inputAll_19_fork_io_outputs_1_rData;
  assign inputAll_20_ready = inputAll_20_fork_io_input_ready;
  always @(*) begin
    inputAll_20_fork_io_outputs_1_ready = inputAll_20_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_20) begin
      inputAll_20_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_20 = (! inputAll_20_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_20_fork_io_outputs_1_m2sPipe_valid = inputAll_20_fork_io_outputs_1_rValid;
  assign inputAll_20_fork_io_outputs_1_m2sPipe_payload = inputAll_20_fork_io_outputs_1_rData;
  assign inputAll_21_ready = inputAll_21_fork_io_input_ready;
  always @(*) begin
    inputAll_21_fork_io_outputs_1_ready = inputAll_21_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_21) begin
      inputAll_21_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_21 = (! inputAll_21_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_21_fork_io_outputs_1_m2sPipe_valid = inputAll_21_fork_io_outputs_1_rValid;
  assign inputAll_21_fork_io_outputs_1_m2sPipe_payload = inputAll_21_fork_io_outputs_1_rData;
  assign inputAll_22_ready = inputAll_22_fork_io_input_ready;
  always @(*) begin
    inputAll_22_fork_io_outputs_1_ready = inputAll_22_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_22) begin
      inputAll_22_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_22 = (! inputAll_22_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_22_fork_io_outputs_1_m2sPipe_valid = inputAll_22_fork_io_outputs_1_rValid;
  assign inputAll_22_fork_io_outputs_1_m2sPipe_payload = inputAll_22_fork_io_outputs_1_rData;
  assign inputAll_23_ready = inputAll_23_fork_io_input_ready;
  always @(*) begin
    inputAll_23_fork_io_outputs_1_ready = inputAll_23_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_23) begin
      inputAll_23_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_23 = (! inputAll_23_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_23_fork_io_outputs_1_m2sPipe_valid = inputAll_23_fork_io_outputs_1_rValid;
  assign inputAll_23_fork_io_outputs_1_m2sPipe_payload = inputAll_23_fork_io_outputs_1_rData;
  assign inputAll_24_ready = inputAll_24_fork_io_input_ready;
  always @(*) begin
    inputAll_24_fork_io_outputs_1_ready = inputAll_24_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_24) begin
      inputAll_24_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_24 = (! inputAll_24_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_24_fork_io_outputs_1_m2sPipe_valid = inputAll_24_fork_io_outputs_1_rValid;
  assign inputAll_24_fork_io_outputs_1_m2sPipe_payload = inputAll_24_fork_io_outputs_1_rData;
  assign inputAll_25_ready = inputAll_25_fork_io_input_ready;
  always @(*) begin
    inputAll_25_fork_io_outputs_1_ready = inputAll_25_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_25) begin
      inputAll_25_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_25 = (! inputAll_25_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_25_fork_io_outputs_1_m2sPipe_valid = inputAll_25_fork_io_outputs_1_rValid;
  assign inputAll_25_fork_io_outputs_1_m2sPipe_payload = inputAll_25_fork_io_outputs_1_rData;
  assign inputAll_26_ready = inputAll_26_fork_io_input_ready;
  always @(*) begin
    inputAll_26_fork_io_outputs_1_ready = inputAll_26_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_26) begin
      inputAll_26_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_26 = (! inputAll_26_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_26_fork_io_outputs_1_m2sPipe_valid = inputAll_26_fork_io_outputs_1_rValid;
  assign inputAll_26_fork_io_outputs_1_m2sPipe_payload = inputAll_26_fork_io_outputs_1_rData;
  assign inputAll_27_ready = inputAll_27_fork_io_input_ready;
  always @(*) begin
    inputAll_27_fork_io_outputs_1_ready = inputAll_27_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_27) begin
      inputAll_27_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_27 = (! inputAll_27_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_27_fork_io_outputs_1_m2sPipe_valid = inputAll_27_fork_io_outputs_1_rValid;
  assign inputAll_27_fork_io_outputs_1_m2sPipe_payload = inputAll_27_fork_io_outputs_1_rData;
  assign inputAll_28_ready = inputAll_28_fork_io_input_ready;
  always @(*) begin
    inputAll_28_fork_io_outputs_1_ready = inputAll_28_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_28) begin
      inputAll_28_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_28 = (! inputAll_28_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_28_fork_io_outputs_1_m2sPipe_valid = inputAll_28_fork_io_outputs_1_rValid;
  assign inputAll_28_fork_io_outputs_1_m2sPipe_payload = inputAll_28_fork_io_outputs_1_rData;
  assign inputAll_29_ready = inputAll_29_fork_io_input_ready;
  always @(*) begin
    inputAll_29_fork_io_outputs_1_ready = inputAll_29_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_29) begin
      inputAll_29_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_29 = (! inputAll_29_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_29_fork_io_outputs_1_m2sPipe_valid = inputAll_29_fork_io_outputs_1_rValid;
  assign inputAll_29_fork_io_outputs_1_m2sPipe_payload = inputAll_29_fork_io_outputs_1_rData;
  assign inputAll_30_ready = inputAll_30_fork_io_input_ready;
  always @(*) begin
    inputAll_30_fork_io_outputs_1_ready = inputAll_30_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_30) begin
      inputAll_30_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_30 = (! inputAll_30_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_30_fork_io_outputs_1_m2sPipe_valid = inputAll_30_fork_io_outputs_1_rValid;
  assign inputAll_30_fork_io_outputs_1_m2sPipe_payload = inputAll_30_fork_io_outputs_1_rData;
  assign inputAll_31_ready = inputAll_31_fork_io_input_ready;
  always @(*) begin
    inputAll_31_fork_io_outputs_1_ready = inputAll_31_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_31) begin
      inputAll_31_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_31 = (! inputAll_31_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_31_fork_io_outputs_1_m2sPipe_valid = inputAll_31_fork_io_outputs_1_rValid;
  assign inputAll_31_fork_io_outputs_1_m2sPipe_payload = inputAll_31_fork_io_outputs_1_rData;
  assign inputAll_32_ready = inputAll_32_fork_io_input_ready;
  always @(*) begin
    inputAll_32_fork_io_outputs_1_ready = inputAll_32_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_32) begin
      inputAll_32_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_32 = (! inputAll_32_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_32_fork_io_outputs_1_m2sPipe_valid = inputAll_32_fork_io_outputs_1_rValid;
  assign inputAll_32_fork_io_outputs_1_m2sPipe_payload = inputAll_32_fork_io_outputs_1_rData;
  assign inputAll_33_ready = inputAll_33_fork_io_input_ready;
  always @(*) begin
    inputAll_33_fork_io_outputs_1_ready = inputAll_33_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_33) begin
      inputAll_33_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_33 = (! inputAll_33_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_33_fork_io_outputs_1_m2sPipe_valid = inputAll_33_fork_io_outputs_1_rValid;
  assign inputAll_33_fork_io_outputs_1_m2sPipe_payload = inputAll_33_fork_io_outputs_1_rData;
  assign inputAll_34_ready = inputAll_34_fork_io_input_ready;
  always @(*) begin
    inputAll_34_fork_io_outputs_1_ready = inputAll_34_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_34) begin
      inputAll_34_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_34 = (! inputAll_34_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_34_fork_io_outputs_1_m2sPipe_valid = inputAll_34_fork_io_outputs_1_rValid;
  assign inputAll_34_fork_io_outputs_1_m2sPipe_payload = inputAll_34_fork_io_outputs_1_rData;
  assign inputAll_35_ready = inputAll_35_fork_io_input_ready;
  always @(*) begin
    inputAll_35_fork_io_outputs_1_ready = inputAll_35_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_35) begin
      inputAll_35_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_35 = (! inputAll_35_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_35_fork_io_outputs_1_m2sPipe_valid = inputAll_35_fork_io_outputs_1_rValid;
  assign inputAll_35_fork_io_outputs_1_m2sPipe_payload = inputAll_35_fork_io_outputs_1_rData;
  assign inputAll_36_ready = inputAll_36_fork_io_input_ready;
  always @(*) begin
    inputAll_36_fork_io_outputs_1_ready = inputAll_36_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_36) begin
      inputAll_36_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_36 = (! inputAll_36_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_36_fork_io_outputs_1_m2sPipe_valid = inputAll_36_fork_io_outputs_1_rValid;
  assign inputAll_36_fork_io_outputs_1_m2sPipe_payload = inputAll_36_fork_io_outputs_1_rData;
  assign inputAll_37_ready = inputAll_37_fork_io_input_ready;
  always @(*) begin
    inputAll_37_fork_io_outputs_1_ready = inputAll_37_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_37) begin
      inputAll_37_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_37 = (! inputAll_37_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_37_fork_io_outputs_1_m2sPipe_valid = inputAll_37_fork_io_outputs_1_rValid;
  assign inputAll_37_fork_io_outputs_1_m2sPipe_payload = inputAll_37_fork_io_outputs_1_rData;
  assign inputAll_38_ready = inputAll_38_fork_io_input_ready;
  always @(*) begin
    inputAll_38_fork_io_outputs_1_ready = inputAll_38_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_38) begin
      inputAll_38_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_38 = (! inputAll_38_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_38_fork_io_outputs_1_m2sPipe_valid = inputAll_38_fork_io_outputs_1_rValid;
  assign inputAll_38_fork_io_outputs_1_m2sPipe_payload = inputAll_38_fork_io_outputs_1_rData;
  assign inputAll_39_ready = inputAll_39_fork_io_input_ready;
  always @(*) begin
    inputAll_39_fork_io_outputs_1_ready = inputAll_39_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_39) begin
      inputAll_39_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_39 = (! inputAll_39_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_39_fork_io_outputs_1_m2sPipe_valid = inputAll_39_fork_io_outputs_1_rValid;
  assign inputAll_39_fork_io_outputs_1_m2sPipe_payload = inputAll_39_fork_io_outputs_1_rData;
  assign inputAll_40_ready = inputAll_40_fork_io_input_ready;
  always @(*) begin
    inputAll_40_fork_io_outputs_1_ready = inputAll_40_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_40) begin
      inputAll_40_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_40 = (! inputAll_40_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_40_fork_io_outputs_1_m2sPipe_valid = inputAll_40_fork_io_outputs_1_rValid;
  assign inputAll_40_fork_io_outputs_1_m2sPipe_payload = inputAll_40_fork_io_outputs_1_rData;
  assign inputAll_41_ready = inputAll_41_fork_io_input_ready;
  always @(*) begin
    inputAll_41_fork_io_outputs_1_ready = inputAll_41_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_41) begin
      inputAll_41_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_41 = (! inputAll_41_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_41_fork_io_outputs_1_m2sPipe_valid = inputAll_41_fork_io_outputs_1_rValid;
  assign inputAll_41_fork_io_outputs_1_m2sPipe_payload = inputAll_41_fork_io_outputs_1_rData;
  assign inputAll_42_ready = inputAll_42_fork_io_input_ready;
  always @(*) begin
    inputAll_42_fork_io_outputs_1_ready = inputAll_42_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_42) begin
      inputAll_42_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_42 = (! inputAll_42_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_42_fork_io_outputs_1_m2sPipe_valid = inputAll_42_fork_io_outputs_1_rValid;
  assign inputAll_42_fork_io_outputs_1_m2sPipe_payload = inputAll_42_fork_io_outputs_1_rData;
  assign inputAll_43_ready = inputAll_43_fork_io_input_ready;
  always @(*) begin
    inputAll_43_fork_io_outputs_1_ready = inputAll_43_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_43) begin
      inputAll_43_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_43 = (! inputAll_43_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_43_fork_io_outputs_1_m2sPipe_valid = inputAll_43_fork_io_outputs_1_rValid;
  assign inputAll_43_fork_io_outputs_1_m2sPipe_payload = inputAll_43_fork_io_outputs_1_rData;
  assign inputAll_44_ready = inputAll_44_fork_io_input_ready;
  always @(*) begin
    inputAll_44_fork_io_outputs_1_ready = inputAll_44_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_44) begin
      inputAll_44_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_44 = (! inputAll_44_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_44_fork_io_outputs_1_m2sPipe_valid = inputAll_44_fork_io_outputs_1_rValid;
  assign inputAll_44_fork_io_outputs_1_m2sPipe_payload = inputAll_44_fork_io_outputs_1_rData;
  assign inputAll_45_ready = inputAll_45_fork_io_input_ready;
  always @(*) begin
    inputAll_45_fork_io_outputs_1_ready = inputAll_45_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_45) begin
      inputAll_45_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_45 = (! inputAll_45_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_45_fork_io_outputs_1_m2sPipe_valid = inputAll_45_fork_io_outputs_1_rValid;
  assign inputAll_45_fork_io_outputs_1_m2sPipe_payload = inputAll_45_fork_io_outputs_1_rData;
  assign inputAll_46_ready = inputAll_46_fork_io_input_ready;
  always @(*) begin
    inputAll_46_fork_io_outputs_1_ready = inputAll_46_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_46) begin
      inputAll_46_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_46 = (! inputAll_46_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_46_fork_io_outputs_1_m2sPipe_valid = inputAll_46_fork_io_outputs_1_rValid;
  assign inputAll_46_fork_io_outputs_1_m2sPipe_payload = inputAll_46_fork_io_outputs_1_rData;
  assign inputAll_47_ready = inputAll_47_fork_io_input_ready;
  always @(*) begin
    inputAll_47_fork_io_outputs_1_ready = inputAll_47_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_47) begin
      inputAll_47_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_47 = (! inputAll_47_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_47_fork_io_outputs_1_m2sPipe_valid = inputAll_47_fork_io_outputs_1_rValid;
  assign inputAll_47_fork_io_outputs_1_m2sPipe_payload = inputAll_47_fork_io_outputs_1_rData;
  assign inputAll_48_ready = inputAll_48_fork_io_input_ready;
  always @(*) begin
    inputAll_48_fork_io_outputs_1_ready = inputAll_48_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_48) begin
      inputAll_48_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_48 = (! inputAll_48_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_48_fork_io_outputs_1_m2sPipe_valid = inputAll_48_fork_io_outputs_1_rValid;
  assign inputAll_48_fork_io_outputs_1_m2sPipe_payload = inputAll_48_fork_io_outputs_1_rData;
  assign inputAll_49_ready = inputAll_49_fork_io_input_ready;
  always @(*) begin
    inputAll_49_fork_io_outputs_1_ready = inputAll_49_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_49) begin
      inputAll_49_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_49 = (! inputAll_49_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_49_fork_io_outputs_1_m2sPipe_valid = inputAll_49_fork_io_outputs_1_rValid;
  assign inputAll_49_fork_io_outputs_1_m2sPipe_payload = inputAll_49_fork_io_outputs_1_rData;
  assign inputAll_50_ready = inputAll_50_fork_io_input_ready;
  always @(*) begin
    inputAll_50_fork_io_outputs_1_ready = inputAll_50_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_50) begin
      inputAll_50_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_50 = (! inputAll_50_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_50_fork_io_outputs_1_m2sPipe_valid = inputAll_50_fork_io_outputs_1_rValid;
  assign inputAll_50_fork_io_outputs_1_m2sPipe_payload = inputAll_50_fork_io_outputs_1_rData;
  assign inputAll_51_ready = inputAll_51_fork_io_input_ready;
  always @(*) begin
    inputAll_51_fork_io_outputs_1_ready = inputAll_51_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_51) begin
      inputAll_51_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_51 = (! inputAll_51_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_51_fork_io_outputs_1_m2sPipe_valid = inputAll_51_fork_io_outputs_1_rValid;
  assign inputAll_51_fork_io_outputs_1_m2sPipe_payload = inputAll_51_fork_io_outputs_1_rData;
  assign inputAll_52_ready = inputAll_52_fork_io_input_ready;
  always @(*) begin
    inputAll_52_fork_io_outputs_1_ready = inputAll_52_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_52) begin
      inputAll_52_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_52 = (! inputAll_52_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_52_fork_io_outputs_1_m2sPipe_valid = inputAll_52_fork_io_outputs_1_rValid;
  assign inputAll_52_fork_io_outputs_1_m2sPipe_payload = inputAll_52_fork_io_outputs_1_rData;
  assign inputAll_53_ready = inputAll_53_fork_io_input_ready;
  always @(*) begin
    inputAll_53_fork_io_outputs_1_ready = inputAll_53_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_53) begin
      inputAll_53_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_53 = (! inputAll_53_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_53_fork_io_outputs_1_m2sPipe_valid = inputAll_53_fork_io_outputs_1_rValid;
  assign inputAll_53_fork_io_outputs_1_m2sPipe_payload = inputAll_53_fork_io_outputs_1_rData;
  assign inputAll_54_ready = inputAll_54_fork_io_input_ready;
  always @(*) begin
    inputAll_54_fork_io_outputs_1_ready = inputAll_54_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_54) begin
      inputAll_54_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_54 = (! inputAll_54_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_54_fork_io_outputs_1_m2sPipe_valid = inputAll_54_fork_io_outputs_1_rValid;
  assign inputAll_54_fork_io_outputs_1_m2sPipe_payload = inputAll_54_fork_io_outputs_1_rData;
  assign inputAll_55_ready = inputAll_55_fork_io_input_ready;
  always @(*) begin
    inputAll_55_fork_io_outputs_1_ready = inputAll_55_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_55) begin
      inputAll_55_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_55 = (! inputAll_55_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_55_fork_io_outputs_1_m2sPipe_valid = inputAll_55_fork_io_outputs_1_rValid;
  assign inputAll_55_fork_io_outputs_1_m2sPipe_payload = inputAll_55_fork_io_outputs_1_rData;
  assign inputAll_56_ready = inputAll_56_fork_io_input_ready;
  always @(*) begin
    inputAll_56_fork_io_outputs_1_ready = inputAll_56_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_56) begin
      inputAll_56_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_56 = (! inputAll_56_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_56_fork_io_outputs_1_m2sPipe_valid = inputAll_56_fork_io_outputs_1_rValid;
  assign inputAll_56_fork_io_outputs_1_m2sPipe_payload = inputAll_56_fork_io_outputs_1_rData;
  assign inputAll_57_ready = inputAll_57_fork_io_input_ready;
  always @(*) begin
    inputAll_57_fork_io_outputs_1_ready = inputAll_57_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_57) begin
      inputAll_57_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_57 = (! inputAll_57_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_57_fork_io_outputs_1_m2sPipe_valid = inputAll_57_fork_io_outputs_1_rValid;
  assign inputAll_57_fork_io_outputs_1_m2sPipe_payload = inputAll_57_fork_io_outputs_1_rData;
  assign inputAll_58_ready = inputAll_58_fork_io_input_ready;
  always @(*) begin
    inputAll_58_fork_io_outputs_1_ready = inputAll_58_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_58) begin
      inputAll_58_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_58 = (! inputAll_58_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_58_fork_io_outputs_1_m2sPipe_valid = inputAll_58_fork_io_outputs_1_rValid;
  assign inputAll_58_fork_io_outputs_1_m2sPipe_payload = inputAll_58_fork_io_outputs_1_rData;
  assign inputAll_59_ready = inputAll_59_fork_io_input_ready;
  always @(*) begin
    inputAll_59_fork_io_outputs_1_ready = inputAll_59_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_59) begin
      inputAll_59_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_59 = (! inputAll_59_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_59_fork_io_outputs_1_m2sPipe_valid = inputAll_59_fork_io_outputs_1_rValid;
  assign inputAll_59_fork_io_outputs_1_m2sPipe_payload = inputAll_59_fork_io_outputs_1_rData;
  assign inputAll_60_ready = inputAll_60_fork_io_input_ready;
  always @(*) begin
    inputAll_60_fork_io_outputs_1_ready = inputAll_60_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_60) begin
      inputAll_60_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_60 = (! inputAll_60_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_60_fork_io_outputs_1_m2sPipe_valid = inputAll_60_fork_io_outputs_1_rValid;
  assign inputAll_60_fork_io_outputs_1_m2sPipe_payload = inputAll_60_fork_io_outputs_1_rData;
  assign inputAll_61_ready = inputAll_61_fork_io_input_ready;
  always @(*) begin
    inputAll_61_fork_io_outputs_1_ready = inputAll_61_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_61) begin
      inputAll_61_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_61 = (! inputAll_61_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_61_fork_io_outputs_1_m2sPipe_valid = inputAll_61_fork_io_outputs_1_rValid;
  assign inputAll_61_fork_io_outputs_1_m2sPipe_payload = inputAll_61_fork_io_outputs_1_rData;
  assign inputAll_62_ready = inputAll_62_fork_io_input_ready;
  always @(*) begin
    inputAll_62_fork_io_outputs_1_ready = inputAll_62_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_62) begin
      inputAll_62_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_62 = (! inputAll_62_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_62_fork_io_outputs_1_m2sPipe_valid = inputAll_62_fork_io_outputs_1_rValid;
  assign inputAll_62_fork_io_outputs_1_m2sPipe_payload = inputAll_62_fork_io_outputs_1_rData;
  assign inputAll_63_ready = inputAll_63_fork_io_input_ready;
  always @(*) begin
    inputAll_63_fork_io_outputs_1_ready = inputAll_63_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_63) begin
      inputAll_63_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_63 = (! inputAll_63_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_63_fork_io_outputs_1_m2sPipe_valid = inputAll_63_fork_io_outputs_1_rValid;
  assign inputAll_63_fork_io_outputs_1_m2sPipe_payload = inputAll_63_fork_io_outputs_1_rData;
  assign inputAll_64_ready = inputAll_64_fork_io_input_ready;
  always @(*) begin
    inputAll_64_fork_io_outputs_1_ready = inputAll_64_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_64) begin
      inputAll_64_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_64 = (! inputAll_64_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_64_fork_io_outputs_1_m2sPipe_valid = inputAll_64_fork_io_outputs_1_rValid;
  assign inputAll_64_fork_io_outputs_1_m2sPipe_payload = inputAll_64_fork_io_outputs_1_rData;
  assign inputAll_65_ready = inputAll_65_fork_io_input_ready;
  always @(*) begin
    inputAll_65_fork_io_outputs_1_ready = inputAll_65_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_65) begin
      inputAll_65_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_65 = (! inputAll_65_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_65_fork_io_outputs_1_m2sPipe_valid = inputAll_65_fork_io_outputs_1_rValid;
  assign inputAll_65_fork_io_outputs_1_m2sPipe_payload = inputAll_65_fork_io_outputs_1_rData;
  assign inputAll_66_ready = inputAll_66_fork_io_input_ready;
  always @(*) begin
    inputAll_66_fork_io_outputs_1_ready = inputAll_66_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_66) begin
      inputAll_66_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_66 = (! inputAll_66_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_66_fork_io_outputs_1_m2sPipe_valid = inputAll_66_fork_io_outputs_1_rValid;
  assign inputAll_66_fork_io_outputs_1_m2sPipe_payload = inputAll_66_fork_io_outputs_1_rData;
  assign inputAll_67_ready = inputAll_67_fork_io_input_ready;
  always @(*) begin
    inputAll_67_fork_io_outputs_1_ready = inputAll_67_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_67) begin
      inputAll_67_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_67 = (! inputAll_67_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_67_fork_io_outputs_1_m2sPipe_valid = inputAll_67_fork_io_outputs_1_rValid;
  assign inputAll_67_fork_io_outputs_1_m2sPipe_payload = inputAll_67_fork_io_outputs_1_rData;
  assign inputAll_68_ready = inputAll_68_fork_io_input_ready;
  always @(*) begin
    inputAll_68_fork_io_outputs_1_ready = inputAll_68_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_68) begin
      inputAll_68_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_68 = (! inputAll_68_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_68_fork_io_outputs_1_m2sPipe_valid = inputAll_68_fork_io_outputs_1_rValid;
  assign inputAll_68_fork_io_outputs_1_m2sPipe_payload = inputAll_68_fork_io_outputs_1_rData;
  assign inputAll_69_ready = inputAll_69_fork_io_input_ready;
  always @(*) begin
    inputAll_69_fork_io_outputs_1_ready = inputAll_69_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_69) begin
      inputAll_69_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_69 = (! inputAll_69_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_69_fork_io_outputs_1_m2sPipe_valid = inputAll_69_fork_io_outputs_1_rValid;
  assign inputAll_69_fork_io_outputs_1_m2sPipe_payload = inputAll_69_fork_io_outputs_1_rData;
  assign inputAll_70_ready = inputAll_70_fork_io_input_ready;
  always @(*) begin
    inputAll_70_fork_io_outputs_1_ready = inputAll_70_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_70) begin
      inputAll_70_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_70 = (! inputAll_70_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_70_fork_io_outputs_1_m2sPipe_valid = inputAll_70_fork_io_outputs_1_rValid;
  assign inputAll_70_fork_io_outputs_1_m2sPipe_payload = inputAll_70_fork_io_outputs_1_rData;
  assign inputAll_71_ready = inputAll_71_fork_io_input_ready;
  always @(*) begin
    inputAll_71_fork_io_outputs_1_ready = inputAll_71_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_71) begin
      inputAll_71_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_71 = (! inputAll_71_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_71_fork_io_outputs_1_m2sPipe_valid = inputAll_71_fork_io_outputs_1_rValid;
  assign inputAll_71_fork_io_outputs_1_m2sPipe_payload = inputAll_71_fork_io_outputs_1_rData;
  assign inputAll_72_ready = inputAll_72_fork_io_input_ready;
  always @(*) begin
    inputAll_72_fork_io_outputs_1_ready = inputAll_72_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_72) begin
      inputAll_72_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_72 = (! inputAll_72_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_72_fork_io_outputs_1_m2sPipe_valid = inputAll_72_fork_io_outputs_1_rValid;
  assign inputAll_72_fork_io_outputs_1_m2sPipe_payload = inputAll_72_fork_io_outputs_1_rData;
  assign inputAll_73_ready = inputAll_73_fork_io_input_ready;
  always @(*) begin
    inputAll_73_fork_io_outputs_1_ready = inputAll_73_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_73) begin
      inputAll_73_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_73 = (! inputAll_73_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_73_fork_io_outputs_1_m2sPipe_valid = inputAll_73_fork_io_outputs_1_rValid;
  assign inputAll_73_fork_io_outputs_1_m2sPipe_payload = inputAll_73_fork_io_outputs_1_rData;
  assign inputAll_74_ready = inputAll_74_fork_io_input_ready;
  always @(*) begin
    inputAll_74_fork_io_outputs_1_ready = inputAll_74_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_74) begin
      inputAll_74_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_74 = (! inputAll_74_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_74_fork_io_outputs_1_m2sPipe_valid = inputAll_74_fork_io_outputs_1_rValid;
  assign inputAll_74_fork_io_outputs_1_m2sPipe_payload = inputAll_74_fork_io_outputs_1_rData;
  assign inputAll_75_ready = inputAll_75_fork_io_input_ready;
  always @(*) begin
    inputAll_75_fork_io_outputs_1_ready = inputAll_75_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_75) begin
      inputAll_75_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_75 = (! inputAll_75_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_75_fork_io_outputs_1_m2sPipe_valid = inputAll_75_fork_io_outputs_1_rValid;
  assign inputAll_75_fork_io_outputs_1_m2sPipe_payload = inputAll_75_fork_io_outputs_1_rData;
  assign inputAll_76_ready = inputAll_76_fork_io_input_ready;
  always @(*) begin
    inputAll_76_fork_io_outputs_1_ready = inputAll_76_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_76) begin
      inputAll_76_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_76 = (! inputAll_76_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_76_fork_io_outputs_1_m2sPipe_valid = inputAll_76_fork_io_outputs_1_rValid;
  assign inputAll_76_fork_io_outputs_1_m2sPipe_payload = inputAll_76_fork_io_outputs_1_rData;
  assign inputAll_77_ready = inputAll_77_fork_io_input_ready;
  always @(*) begin
    inputAll_77_fork_io_outputs_1_ready = inputAll_77_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_77) begin
      inputAll_77_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_77 = (! inputAll_77_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_77_fork_io_outputs_1_m2sPipe_valid = inputAll_77_fork_io_outputs_1_rValid;
  assign inputAll_77_fork_io_outputs_1_m2sPipe_payload = inputAll_77_fork_io_outputs_1_rData;
  assign inputAll_78_ready = inputAll_78_fork_io_input_ready;
  always @(*) begin
    inputAll_78_fork_io_outputs_1_ready = inputAll_78_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_78) begin
      inputAll_78_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_78 = (! inputAll_78_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_78_fork_io_outputs_1_m2sPipe_valid = inputAll_78_fork_io_outputs_1_rValid;
  assign inputAll_78_fork_io_outputs_1_m2sPipe_payload = inputAll_78_fork_io_outputs_1_rData;
  assign inputAll_79_ready = inputAll_79_fork_io_input_ready;
  always @(*) begin
    inputAll_79_fork_io_outputs_1_ready = inputAll_79_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_79) begin
      inputAll_79_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_79 = (! inputAll_79_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_79_fork_io_outputs_1_m2sPipe_valid = inputAll_79_fork_io_outputs_1_rValid;
  assign inputAll_79_fork_io_outputs_1_m2sPipe_payload = inputAll_79_fork_io_outputs_1_rData;
  assign inputAll_80_ready = inputAll_80_fork_io_input_ready;
  always @(*) begin
    inputAll_80_fork_io_outputs_1_ready = inputAll_80_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_80) begin
      inputAll_80_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_80 = (! inputAll_80_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_80_fork_io_outputs_1_m2sPipe_valid = inputAll_80_fork_io_outputs_1_rValid;
  assign inputAll_80_fork_io_outputs_1_m2sPipe_payload = inputAll_80_fork_io_outputs_1_rData;
  assign inputAll_81_ready = inputAll_81_fork_io_input_ready;
  always @(*) begin
    inputAll_81_fork_io_outputs_1_ready = inputAll_81_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_81) begin
      inputAll_81_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_81 = (! inputAll_81_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_81_fork_io_outputs_1_m2sPipe_valid = inputAll_81_fork_io_outputs_1_rValid;
  assign inputAll_81_fork_io_outputs_1_m2sPipe_payload = inputAll_81_fork_io_outputs_1_rData;
  assign inputAll_82_ready = inputAll_82_fork_io_input_ready;
  always @(*) begin
    inputAll_82_fork_io_outputs_1_ready = inputAll_82_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_82) begin
      inputAll_82_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_82 = (! inputAll_82_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_82_fork_io_outputs_1_m2sPipe_valid = inputAll_82_fork_io_outputs_1_rValid;
  assign inputAll_82_fork_io_outputs_1_m2sPipe_payload = inputAll_82_fork_io_outputs_1_rData;
  assign inputAll_83_ready = inputAll_83_fork_io_input_ready;
  always @(*) begin
    inputAll_83_fork_io_outputs_1_ready = inputAll_83_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_83) begin
      inputAll_83_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_83 = (! inputAll_83_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_83_fork_io_outputs_1_m2sPipe_valid = inputAll_83_fork_io_outputs_1_rValid;
  assign inputAll_83_fork_io_outputs_1_m2sPipe_payload = inputAll_83_fork_io_outputs_1_rData;
  assign inputAll_84_ready = inputAll_84_fork_io_input_ready;
  always @(*) begin
    inputAll_84_fork_io_outputs_1_ready = inputAll_84_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_84) begin
      inputAll_84_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_84 = (! inputAll_84_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_84_fork_io_outputs_1_m2sPipe_valid = inputAll_84_fork_io_outputs_1_rValid;
  assign inputAll_84_fork_io_outputs_1_m2sPipe_payload = inputAll_84_fork_io_outputs_1_rData;
  assign inputAll_85_ready = inputAll_85_fork_io_input_ready;
  always @(*) begin
    inputAll_85_fork_io_outputs_1_ready = inputAll_85_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_85) begin
      inputAll_85_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_85 = (! inputAll_85_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_85_fork_io_outputs_1_m2sPipe_valid = inputAll_85_fork_io_outputs_1_rValid;
  assign inputAll_85_fork_io_outputs_1_m2sPipe_payload = inputAll_85_fork_io_outputs_1_rData;
  assign inputAll_86_ready = inputAll_86_fork_io_input_ready;
  always @(*) begin
    inputAll_86_fork_io_outputs_1_ready = inputAll_86_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_86) begin
      inputAll_86_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_86 = (! inputAll_86_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_86_fork_io_outputs_1_m2sPipe_valid = inputAll_86_fork_io_outputs_1_rValid;
  assign inputAll_86_fork_io_outputs_1_m2sPipe_payload = inputAll_86_fork_io_outputs_1_rData;
  assign inputAll_87_ready = inputAll_87_fork_io_input_ready;
  always @(*) begin
    inputAll_87_fork_io_outputs_1_ready = inputAll_87_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_87) begin
      inputAll_87_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_87 = (! inputAll_87_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_87_fork_io_outputs_1_m2sPipe_valid = inputAll_87_fork_io_outputs_1_rValid;
  assign inputAll_87_fork_io_outputs_1_m2sPipe_payload = inputAll_87_fork_io_outputs_1_rData;
  assign inputAll_88_ready = inputAll_88_fork_io_input_ready;
  always @(*) begin
    inputAll_88_fork_io_outputs_1_ready = inputAll_88_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_88) begin
      inputAll_88_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_88 = (! inputAll_88_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_88_fork_io_outputs_1_m2sPipe_valid = inputAll_88_fork_io_outputs_1_rValid;
  assign inputAll_88_fork_io_outputs_1_m2sPipe_payload = inputAll_88_fork_io_outputs_1_rData;
  assign inputAll_89_ready = inputAll_89_fork_io_input_ready;
  always @(*) begin
    inputAll_89_fork_io_outputs_1_ready = inputAll_89_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_89) begin
      inputAll_89_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_89 = (! inputAll_89_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_89_fork_io_outputs_1_m2sPipe_valid = inputAll_89_fork_io_outputs_1_rValid;
  assign inputAll_89_fork_io_outputs_1_m2sPipe_payload = inputAll_89_fork_io_outputs_1_rData;
  assign inputAll_90_ready = inputAll_90_fork_io_input_ready;
  always @(*) begin
    inputAll_90_fork_io_outputs_1_ready = inputAll_90_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_90) begin
      inputAll_90_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_90 = (! inputAll_90_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_90_fork_io_outputs_1_m2sPipe_valid = inputAll_90_fork_io_outputs_1_rValid;
  assign inputAll_90_fork_io_outputs_1_m2sPipe_payload = inputAll_90_fork_io_outputs_1_rData;
  assign inputAll_91_ready = inputAll_91_fork_io_input_ready;
  always @(*) begin
    inputAll_91_fork_io_outputs_1_ready = inputAll_91_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_91) begin
      inputAll_91_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_91 = (! inputAll_91_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_91_fork_io_outputs_1_m2sPipe_valid = inputAll_91_fork_io_outputs_1_rValid;
  assign inputAll_91_fork_io_outputs_1_m2sPipe_payload = inputAll_91_fork_io_outputs_1_rData;
  assign inputAll_92_ready = inputAll_92_fork_io_input_ready;
  always @(*) begin
    inputAll_92_fork_io_outputs_1_ready = inputAll_92_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_92) begin
      inputAll_92_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_92 = (! inputAll_92_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_92_fork_io_outputs_1_m2sPipe_valid = inputAll_92_fork_io_outputs_1_rValid;
  assign inputAll_92_fork_io_outputs_1_m2sPipe_payload = inputAll_92_fork_io_outputs_1_rData;
  assign inputAll_93_ready = inputAll_93_fork_io_input_ready;
  always @(*) begin
    inputAll_93_fork_io_outputs_1_ready = inputAll_93_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_93) begin
      inputAll_93_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_93 = (! inputAll_93_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_93_fork_io_outputs_1_m2sPipe_valid = inputAll_93_fork_io_outputs_1_rValid;
  assign inputAll_93_fork_io_outputs_1_m2sPipe_payload = inputAll_93_fork_io_outputs_1_rData;
  assign inputAll_94_ready = inputAll_94_fork_io_input_ready;
  always @(*) begin
    inputAll_94_fork_io_outputs_1_ready = inputAll_94_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_94) begin
      inputAll_94_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_94 = (! inputAll_94_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_94_fork_io_outputs_1_m2sPipe_valid = inputAll_94_fork_io_outputs_1_rValid;
  assign inputAll_94_fork_io_outputs_1_m2sPipe_payload = inputAll_94_fork_io_outputs_1_rData;
  assign inputAll_95_ready = inputAll_95_fork_io_input_ready;
  always @(*) begin
    inputAll_95_fork_io_outputs_1_ready = inputAll_95_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_95) begin
      inputAll_95_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_95 = (! inputAll_95_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_95_fork_io_outputs_1_m2sPipe_valid = inputAll_95_fork_io_outputs_1_rValid;
  assign inputAll_95_fork_io_outputs_1_m2sPipe_payload = inputAll_95_fork_io_outputs_1_rData;
  assign inputAll_96_ready = inputAll_96_fork_io_input_ready;
  always @(*) begin
    inputAll_96_fork_io_outputs_1_ready = inputAll_96_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_96) begin
      inputAll_96_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_96 = (! inputAll_96_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_96_fork_io_outputs_1_m2sPipe_valid = inputAll_96_fork_io_outputs_1_rValid;
  assign inputAll_96_fork_io_outputs_1_m2sPipe_payload = inputAll_96_fork_io_outputs_1_rData;
  assign inputAll_97_ready = inputAll_97_fork_io_input_ready;
  always @(*) begin
    inputAll_97_fork_io_outputs_1_ready = inputAll_97_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_97) begin
      inputAll_97_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_97 = (! inputAll_97_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_97_fork_io_outputs_1_m2sPipe_valid = inputAll_97_fork_io_outputs_1_rValid;
  assign inputAll_97_fork_io_outputs_1_m2sPipe_payload = inputAll_97_fork_io_outputs_1_rData;
  assign inputAll_98_ready = inputAll_98_fork_io_input_ready;
  always @(*) begin
    inputAll_98_fork_io_outputs_1_ready = inputAll_98_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_98) begin
      inputAll_98_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_98 = (! inputAll_98_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_98_fork_io_outputs_1_m2sPipe_valid = inputAll_98_fork_io_outputs_1_rValid;
  assign inputAll_98_fork_io_outputs_1_m2sPipe_payload = inputAll_98_fork_io_outputs_1_rData;
  assign inputAll_99_ready = inputAll_99_fork_io_input_ready;
  always @(*) begin
    inputAll_99_fork_io_outputs_1_ready = inputAll_99_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_99) begin
      inputAll_99_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_99 = (! inputAll_99_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_99_fork_io_outputs_1_m2sPipe_valid = inputAll_99_fork_io_outputs_1_rValid;
  assign inputAll_99_fork_io_outputs_1_m2sPipe_payload = inputAll_99_fork_io_outputs_1_rData;
  assign inputAll_100_ready = inputAll_100_fork_io_input_ready;
  always @(*) begin
    inputAll_100_fork_io_outputs_1_ready = inputAll_100_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_100) begin
      inputAll_100_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_100 = (! inputAll_100_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_100_fork_io_outputs_1_m2sPipe_valid = inputAll_100_fork_io_outputs_1_rValid;
  assign inputAll_100_fork_io_outputs_1_m2sPipe_payload = inputAll_100_fork_io_outputs_1_rData;
  assign inputAll_101_ready = inputAll_101_fork_io_input_ready;
  always @(*) begin
    inputAll_101_fork_io_outputs_1_ready = inputAll_101_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_101) begin
      inputAll_101_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_101 = (! inputAll_101_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_101_fork_io_outputs_1_m2sPipe_valid = inputAll_101_fork_io_outputs_1_rValid;
  assign inputAll_101_fork_io_outputs_1_m2sPipe_payload = inputAll_101_fork_io_outputs_1_rData;
  assign inputAll_102_ready = inputAll_102_fork_io_input_ready;
  always @(*) begin
    inputAll_102_fork_io_outputs_1_ready = inputAll_102_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_102) begin
      inputAll_102_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_102 = (! inputAll_102_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_102_fork_io_outputs_1_m2sPipe_valid = inputAll_102_fork_io_outputs_1_rValid;
  assign inputAll_102_fork_io_outputs_1_m2sPipe_payload = inputAll_102_fork_io_outputs_1_rData;
  assign inputAll_103_ready = inputAll_103_fork_io_input_ready;
  always @(*) begin
    inputAll_103_fork_io_outputs_1_ready = inputAll_103_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_103) begin
      inputAll_103_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_103 = (! inputAll_103_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_103_fork_io_outputs_1_m2sPipe_valid = inputAll_103_fork_io_outputs_1_rValid;
  assign inputAll_103_fork_io_outputs_1_m2sPipe_payload = inputAll_103_fork_io_outputs_1_rData;
  assign inputAll_104_ready = inputAll_104_fork_io_input_ready;
  always @(*) begin
    inputAll_104_fork_io_outputs_1_ready = inputAll_104_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_104) begin
      inputAll_104_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_104 = (! inputAll_104_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_104_fork_io_outputs_1_m2sPipe_valid = inputAll_104_fork_io_outputs_1_rValid;
  assign inputAll_104_fork_io_outputs_1_m2sPipe_payload = inputAll_104_fork_io_outputs_1_rData;
  assign inputAll_105_ready = inputAll_105_fork_io_input_ready;
  always @(*) begin
    inputAll_105_fork_io_outputs_1_ready = inputAll_105_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_105) begin
      inputAll_105_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_105 = (! inputAll_105_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_105_fork_io_outputs_1_m2sPipe_valid = inputAll_105_fork_io_outputs_1_rValid;
  assign inputAll_105_fork_io_outputs_1_m2sPipe_payload = inputAll_105_fork_io_outputs_1_rData;
  assign inputAll_106_ready = inputAll_106_fork_io_input_ready;
  always @(*) begin
    inputAll_106_fork_io_outputs_1_ready = inputAll_106_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_106) begin
      inputAll_106_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_106 = (! inputAll_106_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_106_fork_io_outputs_1_m2sPipe_valid = inputAll_106_fork_io_outputs_1_rValid;
  assign inputAll_106_fork_io_outputs_1_m2sPipe_payload = inputAll_106_fork_io_outputs_1_rData;
  assign inputAll_107_ready = inputAll_107_fork_io_input_ready;
  always @(*) begin
    inputAll_107_fork_io_outputs_1_ready = inputAll_107_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_107) begin
      inputAll_107_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_107 = (! inputAll_107_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_107_fork_io_outputs_1_m2sPipe_valid = inputAll_107_fork_io_outputs_1_rValid;
  assign inputAll_107_fork_io_outputs_1_m2sPipe_payload = inputAll_107_fork_io_outputs_1_rData;
  assign inputAll_108_ready = inputAll_108_fork_io_input_ready;
  always @(*) begin
    inputAll_108_fork_io_outputs_1_ready = inputAll_108_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_108) begin
      inputAll_108_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_108 = (! inputAll_108_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_108_fork_io_outputs_1_m2sPipe_valid = inputAll_108_fork_io_outputs_1_rValid;
  assign inputAll_108_fork_io_outputs_1_m2sPipe_payload = inputAll_108_fork_io_outputs_1_rData;
  assign inputAll_109_ready = inputAll_109_fork_io_input_ready;
  always @(*) begin
    inputAll_109_fork_io_outputs_1_ready = inputAll_109_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_109) begin
      inputAll_109_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_109 = (! inputAll_109_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_109_fork_io_outputs_1_m2sPipe_valid = inputAll_109_fork_io_outputs_1_rValid;
  assign inputAll_109_fork_io_outputs_1_m2sPipe_payload = inputAll_109_fork_io_outputs_1_rData;
  assign inputAll_110_ready = inputAll_110_fork_io_input_ready;
  always @(*) begin
    inputAll_110_fork_io_outputs_1_ready = inputAll_110_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_110) begin
      inputAll_110_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_110 = (! inputAll_110_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_110_fork_io_outputs_1_m2sPipe_valid = inputAll_110_fork_io_outputs_1_rValid;
  assign inputAll_110_fork_io_outputs_1_m2sPipe_payload = inputAll_110_fork_io_outputs_1_rData;
  assign inputAll_111_ready = inputAll_111_fork_io_input_ready;
  always @(*) begin
    inputAll_111_fork_io_outputs_1_ready = inputAll_111_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_111) begin
      inputAll_111_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_111 = (! inputAll_111_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_111_fork_io_outputs_1_m2sPipe_valid = inputAll_111_fork_io_outputs_1_rValid;
  assign inputAll_111_fork_io_outputs_1_m2sPipe_payload = inputAll_111_fork_io_outputs_1_rData;
  assign inputAll_112_ready = inputAll_112_fork_io_input_ready;
  always @(*) begin
    inputAll_112_fork_io_outputs_1_ready = inputAll_112_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_112) begin
      inputAll_112_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_112 = (! inputAll_112_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_112_fork_io_outputs_1_m2sPipe_valid = inputAll_112_fork_io_outputs_1_rValid;
  assign inputAll_112_fork_io_outputs_1_m2sPipe_payload = inputAll_112_fork_io_outputs_1_rData;
  assign inputAll_113_ready = inputAll_113_fork_io_input_ready;
  always @(*) begin
    inputAll_113_fork_io_outputs_1_ready = inputAll_113_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_113) begin
      inputAll_113_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_113 = (! inputAll_113_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_113_fork_io_outputs_1_m2sPipe_valid = inputAll_113_fork_io_outputs_1_rValid;
  assign inputAll_113_fork_io_outputs_1_m2sPipe_payload = inputAll_113_fork_io_outputs_1_rData;
  assign inputAll_114_ready = inputAll_114_fork_io_input_ready;
  always @(*) begin
    inputAll_114_fork_io_outputs_1_ready = inputAll_114_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_114) begin
      inputAll_114_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_114 = (! inputAll_114_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_114_fork_io_outputs_1_m2sPipe_valid = inputAll_114_fork_io_outputs_1_rValid;
  assign inputAll_114_fork_io_outputs_1_m2sPipe_payload = inputAll_114_fork_io_outputs_1_rData;
  assign inputAll_115_ready = inputAll_115_fork_io_input_ready;
  always @(*) begin
    inputAll_115_fork_io_outputs_1_ready = inputAll_115_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_115) begin
      inputAll_115_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_115 = (! inputAll_115_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_115_fork_io_outputs_1_m2sPipe_valid = inputAll_115_fork_io_outputs_1_rValid;
  assign inputAll_115_fork_io_outputs_1_m2sPipe_payload = inputAll_115_fork_io_outputs_1_rData;
  assign inputAll_116_ready = inputAll_116_fork_io_input_ready;
  always @(*) begin
    inputAll_116_fork_io_outputs_1_ready = inputAll_116_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_116) begin
      inputAll_116_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_116 = (! inputAll_116_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_116_fork_io_outputs_1_m2sPipe_valid = inputAll_116_fork_io_outputs_1_rValid;
  assign inputAll_116_fork_io_outputs_1_m2sPipe_payload = inputAll_116_fork_io_outputs_1_rData;
  assign inputAll_117_ready = inputAll_117_fork_io_input_ready;
  always @(*) begin
    inputAll_117_fork_io_outputs_1_ready = inputAll_117_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_117) begin
      inputAll_117_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_117 = (! inputAll_117_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_117_fork_io_outputs_1_m2sPipe_valid = inputAll_117_fork_io_outputs_1_rValid;
  assign inputAll_117_fork_io_outputs_1_m2sPipe_payload = inputAll_117_fork_io_outputs_1_rData;
  assign inputAll_118_ready = inputAll_118_fork_io_input_ready;
  always @(*) begin
    inputAll_118_fork_io_outputs_1_ready = inputAll_118_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_118) begin
      inputAll_118_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_118 = (! inputAll_118_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_118_fork_io_outputs_1_m2sPipe_valid = inputAll_118_fork_io_outputs_1_rValid;
  assign inputAll_118_fork_io_outputs_1_m2sPipe_payload = inputAll_118_fork_io_outputs_1_rData;
  assign inputAll_119_ready = inputAll_119_fork_io_input_ready;
  always @(*) begin
    inputAll_119_fork_io_outputs_1_ready = inputAll_119_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_119) begin
      inputAll_119_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_119 = (! inputAll_119_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_119_fork_io_outputs_1_m2sPipe_valid = inputAll_119_fork_io_outputs_1_rValid;
  assign inputAll_119_fork_io_outputs_1_m2sPipe_payload = inputAll_119_fork_io_outputs_1_rData;
  assign inputAll_120_ready = inputAll_120_fork_io_input_ready;
  always @(*) begin
    inputAll_120_fork_io_outputs_1_ready = inputAll_120_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_120) begin
      inputAll_120_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_120 = (! inputAll_120_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_120_fork_io_outputs_1_m2sPipe_valid = inputAll_120_fork_io_outputs_1_rValid;
  assign inputAll_120_fork_io_outputs_1_m2sPipe_payload = inputAll_120_fork_io_outputs_1_rData;
  assign inputAll_121_ready = inputAll_121_fork_io_input_ready;
  always @(*) begin
    inputAll_121_fork_io_outputs_1_ready = inputAll_121_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_121) begin
      inputAll_121_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_121 = (! inputAll_121_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_121_fork_io_outputs_1_m2sPipe_valid = inputAll_121_fork_io_outputs_1_rValid;
  assign inputAll_121_fork_io_outputs_1_m2sPipe_payload = inputAll_121_fork_io_outputs_1_rData;
  assign inputAll_122_ready = inputAll_122_fork_io_input_ready;
  always @(*) begin
    inputAll_122_fork_io_outputs_1_ready = inputAll_122_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_122) begin
      inputAll_122_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_122 = (! inputAll_122_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_122_fork_io_outputs_1_m2sPipe_valid = inputAll_122_fork_io_outputs_1_rValid;
  assign inputAll_122_fork_io_outputs_1_m2sPipe_payload = inputAll_122_fork_io_outputs_1_rData;
  assign inputAll_123_ready = inputAll_123_fork_io_input_ready;
  always @(*) begin
    inputAll_123_fork_io_outputs_1_ready = inputAll_123_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_123) begin
      inputAll_123_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_123 = (! inputAll_123_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_123_fork_io_outputs_1_m2sPipe_valid = inputAll_123_fork_io_outputs_1_rValid;
  assign inputAll_123_fork_io_outputs_1_m2sPipe_payload = inputAll_123_fork_io_outputs_1_rData;
  assign inputAll_124_ready = inputAll_124_fork_io_input_ready;
  always @(*) begin
    inputAll_124_fork_io_outputs_1_ready = inputAll_124_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_124) begin
      inputAll_124_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_124 = (! inputAll_124_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_124_fork_io_outputs_1_m2sPipe_valid = inputAll_124_fork_io_outputs_1_rValid;
  assign inputAll_124_fork_io_outputs_1_m2sPipe_payload = inputAll_124_fork_io_outputs_1_rData;
  assign inputAll_125_ready = inputAll_125_fork_io_input_ready;
  always @(*) begin
    inputAll_125_fork_io_outputs_1_ready = inputAll_125_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_125) begin
      inputAll_125_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_125 = (! inputAll_125_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_125_fork_io_outputs_1_m2sPipe_valid = inputAll_125_fork_io_outputs_1_rValid;
  assign inputAll_125_fork_io_outputs_1_m2sPipe_payload = inputAll_125_fork_io_outputs_1_rData;
  assign inputAll_126_ready = inputAll_126_fork_io_input_ready;
  always @(*) begin
    inputAll_126_fork_io_outputs_1_ready = inputAll_126_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_126) begin
      inputAll_126_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_126 = (! inputAll_126_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_126_fork_io_outputs_1_m2sPipe_valid = inputAll_126_fork_io_outputs_1_rValid;
  assign inputAll_126_fork_io_outputs_1_m2sPipe_payload = inputAll_126_fork_io_outputs_1_rData;
  assign inputAll_127_ready = inputAll_127_fork_io_input_ready;
  always @(*) begin
    inputAll_127_fork_io_outputs_1_ready = inputAll_127_fork_io_outputs_1_m2sPipe_ready;
    if(when_Stream_l342_127) begin
      inputAll_127_fork_io_outputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_127 = (! inputAll_127_fork_io_outputs_1_m2sPipe_valid);
  assign inputAll_127_fork_io_outputs_1_m2sPipe_valid = inputAll_127_fork_io_outputs_1_rValid;
  assign inputAll_127_fork_io_outputs_1_m2sPipe_payload = inputAll_127_fork_io_outputs_1_rData;
  assign inputAll_0_valid = io_input_valid;
  assign io_input_ready = inputAll_0_ready;
  assign inputAll_0_payload = io_input_payload;
  assign inputAll_1_valid = inputAll_0_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_0_fork_io_outputs_1_m2sPipe_ready = inputAll_1_ready;
  assign inputAll_1_payload = inputAll_0_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_2_valid = inputAll_1_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_1_fork_io_outputs_1_m2sPipe_ready = inputAll_2_ready;
  assign inputAll_2_payload = inputAll_1_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_3_valid = inputAll_2_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_2_fork_io_outputs_1_m2sPipe_ready = inputAll_3_ready;
  assign inputAll_3_payload = inputAll_2_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_4_valid = inputAll_3_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_3_fork_io_outputs_1_m2sPipe_ready = inputAll_4_ready;
  assign inputAll_4_payload = inputAll_3_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_5_valid = inputAll_4_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_4_fork_io_outputs_1_m2sPipe_ready = inputAll_5_ready;
  assign inputAll_5_payload = inputAll_4_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_6_valid = inputAll_5_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_5_fork_io_outputs_1_m2sPipe_ready = inputAll_6_ready;
  assign inputAll_6_payload = inputAll_5_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_7_valid = inputAll_6_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_6_fork_io_outputs_1_m2sPipe_ready = inputAll_7_ready;
  assign inputAll_7_payload = inputAll_6_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_8_valid = inputAll_7_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_7_fork_io_outputs_1_m2sPipe_ready = inputAll_8_ready;
  assign inputAll_8_payload = inputAll_7_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_9_valid = inputAll_8_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_8_fork_io_outputs_1_m2sPipe_ready = inputAll_9_ready;
  assign inputAll_9_payload = inputAll_8_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_10_valid = inputAll_9_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_9_fork_io_outputs_1_m2sPipe_ready = inputAll_10_ready;
  assign inputAll_10_payload = inputAll_9_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_11_valid = inputAll_10_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_10_fork_io_outputs_1_m2sPipe_ready = inputAll_11_ready;
  assign inputAll_11_payload = inputAll_10_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_12_valid = inputAll_11_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_11_fork_io_outputs_1_m2sPipe_ready = inputAll_12_ready;
  assign inputAll_12_payload = inputAll_11_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_13_valid = inputAll_12_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_12_fork_io_outputs_1_m2sPipe_ready = inputAll_13_ready;
  assign inputAll_13_payload = inputAll_12_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_14_valid = inputAll_13_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_13_fork_io_outputs_1_m2sPipe_ready = inputAll_14_ready;
  assign inputAll_14_payload = inputAll_13_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_15_valid = inputAll_14_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_14_fork_io_outputs_1_m2sPipe_ready = inputAll_15_ready;
  assign inputAll_15_payload = inputAll_14_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_16_valid = inputAll_15_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_15_fork_io_outputs_1_m2sPipe_ready = inputAll_16_ready;
  assign inputAll_16_payload = inputAll_15_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_17_valid = inputAll_16_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_16_fork_io_outputs_1_m2sPipe_ready = inputAll_17_ready;
  assign inputAll_17_payload = inputAll_16_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_18_valid = inputAll_17_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_17_fork_io_outputs_1_m2sPipe_ready = inputAll_18_ready;
  assign inputAll_18_payload = inputAll_17_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_19_valid = inputAll_18_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_18_fork_io_outputs_1_m2sPipe_ready = inputAll_19_ready;
  assign inputAll_19_payload = inputAll_18_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_20_valid = inputAll_19_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_19_fork_io_outputs_1_m2sPipe_ready = inputAll_20_ready;
  assign inputAll_20_payload = inputAll_19_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_21_valid = inputAll_20_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_20_fork_io_outputs_1_m2sPipe_ready = inputAll_21_ready;
  assign inputAll_21_payload = inputAll_20_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_22_valid = inputAll_21_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_21_fork_io_outputs_1_m2sPipe_ready = inputAll_22_ready;
  assign inputAll_22_payload = inputAll_21_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_23_valid = inputAll_22_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_22_fork_io_outputs_1_m2sPipe_ready = inputAll_23_ready;
  assign inputAll_23_payload = inputAll_22_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_24_valid = inputAll_23_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_23_fork_io_outputs_1_m2sPipe_ready = inputAll_24_ready;
  assign inputAll_24_payload = inputAll_23_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_25_valid = inputAll_24_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_24_fork_io_outputs_1_m2sPipe_ready = inputAll_25_ready;
  assign inputAll_25_payload = inputAll_24_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_26_valid = inputAll_25_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_25_fork_io_outputs_1_m2sPipe_ready = inputAll_26_ready;
  assign inputAll_26_payload = inputAll_25_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_27_valid = inputAll_26_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_26_fork_io_outputs_1_m2sPipe_ready = inputAll_27_ready;
  assign inputAll_27_payload = inputAll_26_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_28_valid = inputAll_27_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_27_fork_io_outputs_1_m2sPipe_ready = inputAll_28_ready;
  assign inputAll_28_payload = inputAll_27_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_29_valid = inputAll_28_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_28_fork_io_outputs_1_m2sPipe_ready = inputAll_29_ready;
  assign inputAll_29_payload = inputAll_28_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_30_valid = inputAll_29_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_29_fork_io_outputs_1_m2sPipe_ready = inputAll_30_ready;
  assign inputAll_30_payload = inputAll_29_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_31_valid = inputAll_30_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_30_fork_io_outputs_1_m2sPipe_ready = inputAll_31_ready;
  assign inputAll_31_payload = inputAll_30_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_32_valid = inputAll_31_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_31_fork_io_outputs_1_m2sPipe_ready = inputAll_32_ready;
  assign inputAll_32_payload = inputAll_31_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_33_valid = inputAll_32_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_32_fork_io_outputs_1_m2sPipe_ready = inputAll_33_ready;
  assign inputAll_33_payload = inputAll_32_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_34_valid = inputAll_33_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_33_fork_io_outputs_1_m2sPipe_ready = inputAll_34_ready;
  assign inputAll_34_payload = inputAll_33_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_35_valid = inputAll_34_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_34_fork_io_outputs_1_m2sPipe_ready = inputAll_35_ready;
  assign inputAll_35_payload = inputAll_34_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_36_valid = inputAll_35_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_35_fork_io_outputs_1_m2sPipe_ready = inputAll_36_ready;
  assign inputAll_36_payload = inputAll_35_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_37_valid = inputAll_36_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_36_fork_io_outputs_1_m2sPipe_ready = inputAll_37_ready;
  assign inputAll_37_payload = inputAll_36_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_38_valid = inputAll_37_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_37_fork_io_outputs_1_m2sPipe_ready = inputAll_38_ready;
  assign inputAll_38_payload = inputAll_37_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_39_valid = inputAll_38_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_38_fork_io_outputs_1_m2sPipe_ready = inputAll_39_ready;
  assign inputAll_39_payload = inputAll_38_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_40_valid = inputAll_39_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_39_fork_io_outputs_1_m2sPipe_ready = inputAll_40_ready;
  assign inputAll_40_payload = inputAll_39_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_41_valid = inputAll_40_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_40_fork_io_outputs_1_m2sPipe_ready = inputAll_41_ready;
  assign inputAll_41_payload = inputAll_40_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_42_valid = inputAll_41_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_41_fork_io_outputs_1_m2sPipe_ready = inputAll_42_ready;
  assign inputAll_42_payload = inputAll_41_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_43_valid = inputAll_42_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_42_fork_io_outputs_1_m2sPipe_ready = inputAll_43_ready;
  assign inputAll_43_payload = inputAll_42_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_44_valid = inputAll_43_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_43_fork_io_outputs_1_m2sPipe_ready = inputAll_44_ready;
  assign inputAll_44_payload = inputAll_43_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_45_valid = inputAll_44_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_44_fork_io_outputs_1_m2sPipe_ready = inputAll_45_ready;
  assign inputAll_45_payload = inputAll_44_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_46_valid = inputAll_45_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_45_fork_io_outputs_1_m2sPipe_ready = inputAll_46_ready;
  assign inputAll_46_payload = inputAll_45_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_47_valid = inputAll_46_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_46_fork_io_outputs_1_m2sPipe_ready = inputAll_47_ready;
  assign inputAll_47_payload = inputAll_46_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_48_valid = inputAll_47_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_47_fork_io_outputs_1_m2sPipe_ready = inputAll_48_ready;
  assign inputAll_48_payload = inputAll_47_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_49_valid = inputAll_48_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_48_fork_io_outputs_1_m2sPipe_ready = inputAll_49_ready;
  assign inputAll_49_payload = inputAll_48_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_50_valid = inputAll_49_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_49_fork_io_outputs_1_m2sPipe_ready = inputAll_50_ready;
  assign inputAll_50_payload = inputAll_49_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_51_valid = inputAll_50_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_50_fork_io_outputs_1_m2sPipe_ready = inputAll_51_ready;
  assign inputAll_51_payload = inputAll_50_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_52_valid = inputAll_51_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_51_fork_io_outputs_1_m2sPipe_ready = inputAll_52_ready;
  assign inputAll_52_payload = inputAll_51_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_53_valid = inputAll_52_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_52_fork_io_outputs_1_m2sPipe_ready = inputAll_53_ready;
  assign inputAll_53_payload = inputAll_52_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_54_valid = inputAll_53_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_53_fork_io_outputs_1_m2sPipe_ready = inputAll_54_ready;
  assign inputAll_54_payload = inputAll_53_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_55_valid = inputAll_54_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_54_fork_io_outputs_1_m2sPipe_ready = inputAll_55_ready;
  assign inputAll_55_payload = inputAll_54_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_56_valid = inputAll_55_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_55_fork_io_outputs_1_m2sPipe_ready = inputAll_56_ready;
  assign inputAll_56_payload = inputAll_55_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_57_valid = inputAll_56_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_56_fork_io_outputs_1_m2sPipe_ready = inputAll_57_ready;
  assign inputAll_57_payload = inputAll_56_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_58_valid = inputAll_57_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_57_fork_io_outputs_1_m2sPipe_ready = inputAll_58_ready;
  assign inputAll_58_payload = inputAll_57_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_59_valid = inputAll_58_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_58_fork_io_outputs_1_m2sPipe_ready = inputAll_59_ready;
  assign inputAll_59_payload = inputAll_58_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_60_valid = inputAll_59_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_59_fork_io_outputs_1_m2sPipe_ready = inputAll_60_ready;
  assign inputAll_60_payload = inputAll_59_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_61_valid = inputAll_60_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_60_fork_io_outputs_1_m2sPipe_ready = inputAll_61_ready;
  assign inputAll_61_payload = inputAll_60_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_62_valid = inputAll_61_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_61_fork_io_outputs_1_m2sPipe_ready = inputAll_62_ready;
  assign inputAll_62_payload = inputAll_61_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_63_valid = inputAll_62_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_62_fork_io_outputs_1_m2sPipe_ready = inputAll_63_ready;
  assign inputAll_63_payload = inputAll_62_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_64_valid = inputAll_63_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_63_fork_io_outputs_1_m2sPipe_ready = inputAll_64_ready;
  assign inputAll_64_payload = inputAll_63_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_65_valid = inputAll_64_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_64_fork_io_outputs_1_m2sPipe_ready = inputAll_65_ready;
  assign inputAll_65_payload = inputAll_64_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_66_valid = inputAll_65_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_65_fork_io_outputs_1_m2sPipe_ready = inputAll_66_ready;
  assign inputAll_66_payload = inputAll_65_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_67_valid = inputAll_66_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_66_fork_io_outputs_1_m2sPipe_ready = inputAll_67_ready;
  assign inputAll_67_payload = inputAll_66_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_68_valid = inputAll_67_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_67_fork_io_outputs_1_m2sPipe_ready = inputAll_68_ready;
  assign inputAll_68_payload = inputAll_67_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_69_valid = inputAll_68_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_68_fork_io_outputs_1_m2sPipe_ready = inputAll_69_ready;
  assign inputAll_69_payload = inputAll_68_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_70_valid = inputAll_69_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_69_fork_io_outputs_1_m2sPipe_ready = inputAll_70_ready;
  assign inputAll_70_payload = inputAll_69_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_71_valid = inputAll_70_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_70_fork_io_outputs_1_m2sPipe_ready = inputAll_71_ready;
  assign inputAll_71_payload = inputAll_70_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_72_valid = inputAll_71_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_71_fork_io_outputs_1_m2sPipe_ready = inputAll_72_ready;
  assign inputAll_72_payload = inputAll_71_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_73_valid = inputAll_72_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_72_fork_io_outputs_1_m2sPipe_ready = inputAll_73_ready;
  assign inputAll_73_payload = inputAll_72_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_74_valid = inputAll_73_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_73_fork_io_outputs_1_m2sPipe_ready = inputAll_74_ready;
  assign inputAll_74_payload = inputAll_73_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_75_valid = inputAll_74_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_74_fork_io_outputs_1_m2sPipe_ready = inputAll_75_ready;
  assign inputAll_75_payload = inputAll_74_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_76_valid = inputAll_75_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_75_fork_io_outputs_1_m2sPipe_ready = inputAll_76_ready;
  assign inputAll_76_payload = inputAll_75_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_77_valid = inputAll_76_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_76_fork_io_outputs_1_m2sPipe_ready = inputAll_77_ready;
  assign inputAll_77_payload = inputAll_76_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_78_valid = inputAll_77_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_77_fork_io_outputs_1_m2sPipe_ready = inputAll_78_ready;
  assign inputAll_78_payload = inputAll_77_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_79_valid = inputAll_78_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_78_fork_io_outputs_1_m2sPipe_ready = inputAll_79_ready;
  assign inputAll_79_payload = inputAll_78_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_80_valid = inputAll_79_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_79_fork_io_outputs_1_m2sPipe_ready = inputAll_80_ready;
  assign inputAll_80_payload = inputAll_79_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_81_valid = inputAll_80_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_80_fork_io_outputs_1_m2sPipe_ready = inputAll_81_ready;
  assign inputAll_81_payload = inputAll_80_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_82_valid = inputAll_81_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_81_fork_io_outputs_1_m2sPipe_ready = inputAll_82_ready;
  assign inputAll_82_payload = inputAll_81_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_83_valid = inputAll_82_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_82_fork_io_outputs_1_m2sPipe_ready = inputAll_83_ready;
  assign inputAll_83_payload = inputAll_82_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_84_valid = inputAll_83_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_83_fork_io_outputs_1_m2sPipe_ready = inputAll_84_ready;
  assign inputAll_84_payload = inputAll_83_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_85_valid = inputAll_84_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_84_fork_io_outputs_1_m2sPipe_ready = inputAll_85_ready;
  assign inputAll_85_payload = inputAll_84_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_86_valid = inputAll_85_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_85_fork_io_outputs_1_m2sPipe_ready = inputAll_86_ready;
  assign inputAll_86_payload = inputAll_85_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_87_valid = inputAll_86_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_86_fork_io_outputs_1_m2sPipe_ready = inputAll_87_ready;
  assign inputAll_87_payload = inputAll_86_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_88_valid = inputAll_87_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_87_fork_io_outputs_1_m2sPipe_ready = inputAll_88_ready;
  assign inputAll_88_payload = inputAll_87_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_89_valid = inputAll_88_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_88_fork_io_outputs_1_m2sPipe_ready = inputAll_89_ready;
  assign inputAll_89_payload = inputAll_88_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_90_valid = inputAll_89_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_89_fork_io_outputs_1_m2sPipe_ready = inputAll_90_ready;
  assign inputAll_90_payload = inputAll_89_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_91_valid = inputAll_90_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_90_fork_io_outputs_1_m2sPipe_ready = inputAll_91_ready;
  assign inputAll_91_payload = inputAll_90_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_92_valid = inputAll_91_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_91_fork_io_outputs_1_m2sPipe_ready = inputAll_92_ready;
  assign inputAll_92_payload = inputAll_91_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_93_valid = inputAll_92_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_92_fork_io_outputs_1_m2sPipe_ready = inputAll_93_ready;
  assign inputAll_93_payload = inputAll_92_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_94_valid = inputAll_93_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_93_fork_io_outputs_1_m2sPipe_ready = inputAll_94_ready;
  assign inputAll_94_payload = inputAll_93_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_95_valid = inputAll_94_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_94_fork_io_outputs_1_m2sPipe_ready = inputAll_95_ready;
  assign inputAll_95_payload = inputAll_94_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_96_valid = inputAll_95_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_95_fork_io_outputs_1_m2sPipe_ready = inputAll_96_ready;
  assign inputAll_96_payload = inputAll_95_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_97_valid = inputAll_96_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_96_fork_io_outputs_1_m2sPipe_ready = inputAll_97_ready;
  assign inputAll_97_payload = inputAll_96_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_98_valid = inputAll_97_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_97_fork_io_outputs_1_m2sPipe_ready = inputAll_98_ready;
  assign inputAll_98_payload = inputAll_97_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_99_valid = inputAll_98_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_98_fork_io_outputs_1_m2sPipe_ready = inputAll_99_ready;
  assign inputAll_99_payload = inputAll_98_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_100_valid = inputAll_99_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_99_fork_io_outputs_1_m2sPipe_ready = inputAll_100_ready;
  assign inputAll_100_payload = inputAll_99_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_101_valid = inputAll_100_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_100_fork_io_outputs_1_m2sPipe_ready = inputAll_101_ready;
  assign inputAll_101_payload = inputAll_100_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_102_valid = inputAll_101_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_101_fork_io_outputs_1_m2sPipe_ready = inputAll_102_ready;
  assign inputAll_102_payload = inputAll_101_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_103_valid = inputAll_102_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_102_fork_io_outputs_1_m2sPipe_ready = inputAll_103_ready;
  assign inputAll_103_payload = inputAll_102_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_104_valid = inputAll_103_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_103_fork_io_outputs_1_m2sPipe_ready = inputAll_104_ready;
  assign inputAll_104_payload = inputAll_103_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_105_valid = inputAll_104_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_104_fork_io_outputs_1_m2sPipe_ready = inputAll_105_ready;
  assign inputAll_105_payload = inputAll_104_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_106_valid = inputAll_105_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_105_fork_io_outputs_1_m2sPipe_ready = inputAll_106_ready;
  assign inputAll_106_payload = inputAll_105_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_107_valid = inputAll_106_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_106_fork_io_outputs_1_m2sPipe_ready = inputAll_107_ready;
  assign inputAll_107_payload = inputAll_106_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_108_valid = inputAll_107_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_107_fork_io_outputs_1_m2sPipe_ready = inputAll_108_ready;
  assign inputAll_108_payload = inputAll_107_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_109_valid = inputAll_108_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_108_fork_io_outputs_1_m2sPipe_ready = inputAll_109_ready;
  assign inputAll_109_payload = inputAll_108_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_110_valid = inputAll_109_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_109_fork_io_outputs_1_m2sPipe_ready = inputAll_110_ready;
  assign inputAll_110_payload = inputAll_109_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_111_valid = inputAll_110_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_110_fork_io_outputs_1_m2sPipe_ready = inputAll_111_ready;
  assign inputAll_111_payload = inputAll_110_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_112_valid = inputAll_111_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_111_fork_io_outputs_1_m2sPipe_ready = inputAll_112_ready;
  assign inputAll_112_payload = inputAll_111_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_113_valid = inputAll_112_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_112_fork_io_outputs_1_m2sPipe_ready = inputAll_113_ready;
  assign inputAll_113_payload = inputAll_112_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_114_valid = inputAll_113_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_113_fork_io_outputs_1_m2sPipe_ready = inputAll_114_ready;
  assign inputAll_114_payload = inputAll_113_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_115_valid = inputAll_114_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_114_fork_io_outputs_1_m2sPipe_ready = inputAll_115_ready;
  assign inputAll_115_payload = inputAll_114_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_116_valid = inputAll_115_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_115_fork_io_outputs_1_m2sPipe_ready = inputAll_116_ready;
  assign inputAll_116_payload = inputAll_115_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_117_valid = inputAll_116_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_116_fork_io_outputs_1_m2sPipe_ready = inputAll_117_ready;
  assign inputAll_117_payload = inputAll_116_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_118_valid = inputAll_117_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_117_fork_io_outputs_1_m2sPipe_ready = inputAll_118_ready;
  assign inputAll_118_payload = inputAll_117_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_119_valid = inputAll_118_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_118_fork_io_outputs_1_m2sPipe_ready = inputAll_119_ready;
  assign inputAll_119_payload = inputAll_118_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_120_valid = inputAll_119_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_119_fork_io_outputs_1_m2sPipe_ready = inputAll_120_ready;
  assign inputAll_120_payload = inputAll_119_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_121_valid = inputAll_120_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_120_fork_io_outputs_1_m2sPipe_ready = inputAll_121_ready;
  assign inputAll_121_payload = inputAll_120_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_122_valid = inputAll_121_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_121_fork_io_outputs_1_m2sPipe_ready = inputAll_122_ready;
  assign inputAll_122_payload = inputAll_121_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_123_valid = inputAll_122_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_122_fork_io_outputs_1_m2sPipe_ready = inputAll_123_ready;
  assign inputAll_123_payload = inputAll_122_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_124_valid = inputAll_123_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_123_fork_io_outputs_1_m2sPipe_ready = inputAll_124_ready;
  assign inputAll_124_payload = inputAll_123_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_125_valid = inputAll_124_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_124_fork_io_outputs_1_m2sPipe_ready = inputAll_125_ready;
  assign inputAll_125_payload = inputAll_124_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_126_valid = inputAll_125_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_125_fork_io_outputs_1_m2sPipe_ready = inputAll_126_ready;
  assign inputAll_126_payload = inputAll_125_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_127_valid = inputAll_126_fork_io_outputs_1_m2sPipe_valid;
  assign inputAll_126_fork_io_outputs_1_m2sPipe_ready = inputAll_127_ready;
  assign inputAll_127_payload = inputAll_126_fork_io_outputs_1_m2sPipe_payload;
  assign inputAll_127_fork_io_outputs_1_m2sPipe_ready = 1'b1;
  assign mulResGroup_0_valid = (inputAll_0_fork_io_outputs_0_valid && inputAll_127_fork_io_outputs_0_valid);
  assign mulResGroup_0_payload = {{13{_zz_mulResGroup_0_payload[8]}}, _zz_mulResGroup_0_payload};
  assign mulResGroup_1_valid = (inputAll_1_fork_io_outputs_0_valid && inputAll_126_fork_io_outputs_0_valid);
  assign mulResGroup_1_payload = {{13{_zz_mulResGroup_1_payload[8]}}, _zz_mulResGroup_1_payload};
  assign mulResGroup_2_valid = (inputAll_2_fork_io_outputs_0_valid && inputAll_125_fork_io_outputs_0_valid);
  assign mulResGroup_2_payload = {{13{_zz_mulResGroup_2_payload[8]}}, _zz_mulResGroup_2_payload};
  assign mulResGroup_3_valid = (inputAll_3_fork_io_outputs_0_valid && inputAll_124_fork_io_outputs_0_valid);
  assign mulResGroup_3_payload = {{13{_zz_mulResGroup_3_payload[8]}}, _zz_mulResGroup_3_payload};
  assign mulResGroup_4_valid = (inputAll_4_fork_io_outputs_0_valid && inputAll_123_fork_io_outputs_0_valid);
  assign mulResGroup_4_payload = {{13{_zz_mulResGroup_4_payload[8]}}, _zz_mulResGroup_4_payload};
  assign mulResGroup_5_valid = (inputAll_5_fork_io_outputs_0_valid && inputAll_122_fork_io_outputs_0_valid);
  assign mulResGroup_5_payload = {{13{_zz_mulResGroup_5_payload[8]}}, _zz_mulResGroup_5_payload};
  assign mulResGroup_6_valid = (inputAll_6_fork_io_outputs_0_valid && inputAll_121_fork_io_outputs_0_valid);
  assign mulResGroup_6_payload = {{13{_zz_mulResGroup_6_payload[8]}}, _zz_mulResGroup_6_payload};
  assign mulResGroup_7_valid = (inputAll_7_fork_io_outputs_0_valid && inputAll_120_fork_io_outputs_0_valid);
  assign mulResGroup_7_payload = {{13{_zz_mulResGroup_7_payload[8]}}, _zz_mulResGroup_7_payload};
  assign mulResGroup_8_valid = (inputAll_8_fork_io_outputs_0_valid && inputAll_119_fork_io_outputs_0_valid);
  assign mulResGroup_8_payload = {{13{_zz_mulResGroup_8_payload[8]}}, _zz_mulResGroup_8_payload};
  assign mulResGroup_9_valid = (inputAll_9_fork_io_outputs_0_valid && inputAll_118_fork_io_outputs_0_valid);
  assign mulResGroup_9_payload = {{13{_zz_mulResGroup_9_payload[8]}}, _zz_mulResGroup_9_payload};
  assign mulResGroup_10_valid = (inputAll_10_fork_io_outputs_0_valid && inputAll_117_fork_io_outputs_0_valid);
  assign mulResGroup_10_payload = {{13{_zz_mulResGroup_10_payload[8]}}, _zz_mulResGroup_10_payload};
  assign mulResGroup_11_valid = (inputAll_11_fork_io_outputs_0_valid && inputAll_116_fork_io_outputs_0_valid);
  assign mulResGroup_11_payload = {{13{_zz_mulResGroup_11_payload[8]}}, _zz_mulResGroup_11_payload};
  assign mulResGroup_12_valid = (inputAll_12_fork_io_outputs_0_valid && inputAll_115_fork_io_outputs_0_valid);
  assign mulResGroup_12_payload = {{13{_zz_mulResGroup_12_payload[8]}}, _zz_mulResGroup_12_payload};
  assign mulResGroup_13_valid = (inputAll_13_fork_io_outputs_0_valid && inputAll_114_fork_io_outputs_0_valid);
  assign mulResGroup_13_payload = {{13{_zz_mulResGroup_13_payload[8]}}, _zz_mulResGroup_13_payload};
  assign mulResGroup_14_valid = (inputAll_14_fork_io_outputs_0_valid && inputAll_113_fork_io_outputs_0_valid);
  assign mulResGroup_14_payload = {{13{_zz_mulResGroup_14_payload[8]}}, _zz_mulResGroup_14_payload};
  assign mulResGroup_15_valid = (inputAll_15_fork_io_outputs_0_valid && inputAll_112_fork_io_outputs_0_valid);
  assign mulResGroup_15_payload = {{13{_zz_mulResGroup_15_payload[8]}}, _zz_mulResGroup_15_payload};
  assign mulResGroup_16_valid = (inputAll_16_fork_io_outputs_0_valid && inputAll_111_fork_io_outputs_0_valid);
  assign mulResGroup_16_payload = {{12{_zz_mulResGroup_16_payload[9]}}, _zz_mulResGroup_16_payload};
  assign mulResGroup_17_valid = (inputAll_17_fork_io_outputs_0_valid && inputAll_110_fork_io_outputs_0_valid);
  assign mulResGroup_17_payload = {{12{_zz_mulResGroup_17_payload[9]}}, _zz_mulResGroup_17_payload};
  assign mulResGroup_18_valid = (inputAll_18_fork_io_outputs_0_valid && inputAll_109_fork_io_outputs_0_valid);
  assign mulResGroup_18_payload = {{12{_zz_mulResGroup_18_payload[9]}}, _zz_mulResGroup_18_payload};
  assign mulResGroup_19_valid = (inputAll_19_fork_io_outputs_0_valid && inputAll_108_fork_io_outputs_0_valid);
  assign mulResGroup_19_payload = {{13{_zz_mulResGroup_19_payload[8]}}, _zz_mulResGroup_19_payload};
  assign mulResGroup_20_valid = (inputAll_20_fork_io_outputs_0_valid && inputAll_107_fork_io_outputs_0_valid);
  assign mulResGroup_20_payload = {{13{_zz_mulResGroup_20_payload[8]}}, _zz_mulResGroup_20_payload};
  assign mulResGroup_21_valid = (inputAll_21_fork_io_outputs_0_valid && inputAll_106_fork_io_outputs_0_valid);
  assign mulResGroup_21_payload = {{11{_zz_mulResGroup_21_payload[10]}}, _zz_mulResGroup_21_payload};
  assign mulResGroup_22_valid = (inputAll_22_fork_io_outputs_0_valid && inputAll_105_fork_io_outputs_0_valid);
  assign mulResGroup_22_payload = {{11{_zz_mulResGroup_22_payload[10]}}, _zz_mulResGroup_22_payload};
  assign mulResGroup_23_valid = (inputAll_23_fork_io_outputs_0_valid && inputAll_104_fork_io_outputs_0_valid);
  assign mulResGroup_23_payload = {{11{_zz_mulResGroup_23_payload[10]}}, _zz_mulResGroup_23_payload};
  assign mulResGroup_24_valid = (inputAll_24_fork_io_outputs_0_valid && inputAll_103_fork_io_outputs_0_valid);
  assign mulResGroup_24_payload = {{11{_zz_mulResGroup_24_payload[10]}}, _zz_mulResGroup_24_payload};
  assign mulResGroup_25_valid = (inputAll_25_fork_io_outputs_0_valid && inputAll_102_fork_io_outputs_0_valid);
  assign mulResGroup_25_payload = {{11{_zz_mulResGroup_25_payload[10]}}, _zz_mulResGroup_25_payload};
  assign mulResGroup_26_valid = (inputAll_26_fork_io_outputs_0_valid && inputAll_101_fork_io_outputs_0_valid);
  assign mulResGroup_26_payload = {{13{_zz_mulResGroup_26_payload[8]}}, _zz_mulResGroup_26_payload};
  assign mulResGroup_27_valid = (inputAll_27_fork_io_outputs_0_valid && inputAll_100_fork_io_outputs_0_valid);
  assign mulResGroup_27_payload = {{12{_zz_mulResGroup_27_payload[9]}}, _zz_mulResGroup_27_payload};
  assign mulResGroup_28_valid = (inputAll_28_fork_io_outputs_0_valid && inputAll_99_fork_io_outputs_0_valid);
  assign mulResGroup_28_payload = {{11{_zz_mulResGroup_28_payload[10]}}, _zz_mulResGroup_28_payload};
  assign mulResGroup_29_valid = (inputAll_29_fork_io_outputs_0_valid && inputAll_98_fork_io_outputs_0_valid);
  assign mulResGroup_29_payload = {{11{_zz_mulResGroup_29_payload[10]}}, _zz_mulResGroup_29_payload};
  assign mulResGroup_30_valid = (inputAll_30_fork_io_outputs_0_valid && inputAll_97_fork_io_outputs_0_valid);
  assign mulResGroup_30_payload = {{11{_zz_mulResGroup_30_payload[10]}}, _zz_mulResGroup_30_payload};
  assign mulResGroup_31_valid = (inputAll_31_fork_io_outputs_0_valid && inputAll_96_fork_io_outputs_0_valid);
  assign mulResGroup_31_payload = {{11{_zz_mulResGroup_31_payload[10]}}, _zz_mulResGroup_31_payload};
  assign mulResGroup_32_valid = (inputAll_32_fork_io_outputs_0_valid && inputAll_95_fork_io_outputs_0_valid);
  assign mulResGroup_32_payload = {{13{_zz_mulResGroup_32_payload[8]}}, _zz_mulResGroup_32_payload};
  assign mulResGroup_33_valid = (inputAll_33_fork_io_outputs_0_valid && inputAll_94_fork_io_outputs_0_valid);
  assign mulResGroup_33_payload = {{11{_zz_mulResGroup_33_payload[10]}}, _zz_mulResGroup_33_payload};
  assign mulResGroup_34_valid = (inputAll_34_fork_io_outputs_0_valid && inputAll_93_fork_io_outputs_0_valid);
  assign mulResGroup_34_payload = {{10{_zz_mulResGroup_34_payload[11]}}, _zz_mulResGroup_34_payload};
  assign mulResGroup_35_valid = (inputAll_35_fork_io_outputs_0_valid && inputAll_92_fork_io_outputs_0_valid);
  assign mulResGroup_35_payload = {{10{_zz_mulResGroup_35_payload[11]}}, _zz_mulResGroup_35_payload};
  assign mulResGroup_36_valid = (inputAll_36_fork_io_outputs_0_valid && inputAll_91_fork_io_outputs_0_valid);
  assign mulResGroup_36_payload = {{9{_zz_mulResGroup_36_payload[12]}}, _zz_mulResGroup_36_payload};
  assign mulResGroup_37_valid = (inputAll_37_fork_io_outputs_0_valid && inputAll_90_fork_io_outputs_0_valid);
  assign mulResGroup_37_payload = {{10{_zz_mulResGroup_37_payload[11]}}, _zz_mulResGroup_37_payload};
  assign mulResGroup_38_valid = (inputAll_38_fork_io_outputs_0_valid && inputAll_89_fork_io_outputs_0_valid);
  assign mulResGroup_38_payload = {{11{_zz_mulResGroup_38_payload[10]}}, _zz_mulResGroup_38_payload};
  assign mulResGroup_39_valid = (inputAll_39_fork_io_outputs_0_valid && inputAll_88_fork_io_outputs_0_valid);
  assign mulResGroup_39_payload = {{12{_zz_mulResGroup_39_payload[9]}}, _zz_mulResGroup_39_payload};
  assign mulResGroup_40_valid = (inputAll_40_fork_io_outputs_0_valid && inputAll_87_fork_io_outputs_0_valid);
  assign mulResGroup_40_payload = {{10{_zz_mulResGroup_40_payload[11]}}, _zz_mulResGroup_40_payload};
  assign mulResGroup_41_valid = (inputAll_41_fork_io_outputs_0_valid && inputAll_86_fork_io_outputs_0_valid);
  assign mulResGroup_41_payload = {{9{_zz_mulResGroup_41_payload[12]}}, _zz_mulResGroup_41_payload};
  assign mulResGroup_42_valid = (inputAll_42_fork_io_outputs_0_valid && inputAll_85_fork_io_outputs_0_valid);
  assign mulResGroup_42_payload = {{9{_zz_mulResGroup_42_payload[12]}}, _zz_mulResGroup_42_payload};
  assign mulResGroup_43_valid = (inputAll_43_fork_io_outputs_0_valid && inputAll_84_fork_io_outputs_0_valid);
  assign mulResGroup_43_payload = {{9{_zz_mulResGroup_43_payload[12]}}, _zz_mulResGroup_43_payload};
  assign mulResGroup_44_valid = (inputAll_44_fork_io_outputs_0_valid && inputAll_83_fork_io_outputs_0_valid);
  assign mulResGroup_44_payload = {{11{_zz_mulResGroup_44_payload[10]}}, _zz_mulResGroup_44_payload};
  assign mulResGroup_45_valid = (inputAll_45_fork_io_outputs_0_valid && inputAll_82_fork_io_outputs_0_valid);
  assign mulResGroup_45_payload = {{11{_zz_mulResGroup_45_payload[10]}}, _zz_mulResGroup_45_payload};
  assign mulResGroup_46_valid = (inputAll_46_fork_io_outputs_0_valid && inputAll_81_fork_io_outputs_0_valid);
  assign mulResGroup_46_payload = {{9{_zz_mulResGroup_46_payload[12]}}, _zz_mulResGroup_46_payload};
  assign mulResGroup_47_valid = (inputAll_47_fork_io_outputs_0_valid && inputAll_80_fork_io_outputs_0_valid);
  assign mulResGroup_47_payload = {{8{_zz_mulResGroup_47_payload[13]}}, _zz_mulResGroup_47_payload};
  assign mulResGroup_48_valid = (inputAll_48_fork_io_outputs_0_valid && inputAll_79_fork_io_outputs_0_valid);
  assign mulResGroup_48_payload = {{8{_zz_mulResGroup_48_payload[13]}}, _zz_mulResGroup_48_payload};
  assign mulResGroup_49_valid = (inputAll_49_fork_io_outputs_0_valid && inputAll_78_fork_io_outputs_0_valid);
  assign mulResGroup_49_payload = {{8{_zz_mulResGroup_49_payload[13]}}, _zz_mulResGroup_49_payload};
  assign mulResGroup_50_valid = (inputAll_50_fork_io_outputs_0_valid && inputAll_77_fork_io_outputs_0_valid);
  assign mulResGroup_50_payload = {{9{_zz_mulResGroup_50_payload[12]}}, _zz_mulResGroup_50_payload};
  assign mulResGroup_51_valid = (inputAll_51_fork_io_outputs_0_valid && inputAll_76_fork_io_outputs_0_valid);
  assign mulResGroup_51_payload = {{13{_zz_mulResGroup_51_payload[8]}}, _zz_mulResGroup_51_payload};
  assign mulResGroup_52_valid = (inputAll_52_fork_io_outputs_0_valid && inputAll_75_fork_io_outputs_0_valid);
  assign mulResGroup_52_payload = {{9{_zz_mulResGroup_52_payload[12]}}, _zz_mulResGroup_52_payload};
  assign mulResGroup_53_valid = (inputAll_53_fork_io_outputs_0_valid && inputAll_74_fork_io_outputs_0_valid);
  assign mulResGroup_53_payload = {{8{_zz_mulResGroup_53_payload[13]}}, _zz_mulResGroup_53_payload};
  assign mulResGroup_54_valid = (inputAll_54_fork_io_outputs_0_valid && inputAll_73_fork_io_outputs_0_valid);
  assign mulResGroup_54_payload = {{8{_zz_mulResGroup_54_payload[13]}}, _zz_mulResGroup_54_payload};
  assign mulResGroup_55_valid = (inputAll_55_fork_io_outputs_0_valid && inputAll_72_fork_io_outputs_0_valid);
  assign mulResGroup_55_payload = {{7{_zz_mulResGroup_55_payload[14]}}, _zz_mulResGroup_55_payload};
  assign mulResGroup_56_valid = (inputAll_56_fork_io_outputs_0_valid && inputAll_71_fork_io_outputs_0_valid);
  assign mulResGroup_56_payload = {{8{_zz_mulResGroup_56_payload[13]}}, _zz_mulResGroup_56_payload};
  assign mulResGroup_57_valid = (inputAll_57_fork_io_outputs_0_valid && inputAll_70_fork_io_outputs_0_valid);
  assign mulResGroup_57_payload = {{10{_zz_mulResGroup_57_payload[11]}}, _zz_mulResGroup_57_payload};
  assign mulResGroup_58_valid = (inputAll_58_fork_io_outputs_0_valid && inputAll_69_fork_io_outputs_0_valid);
  assign mulResGroup_58_payload = {{8{_zz_mulResGroup_58_payload[13]}}, _zz_mulResGroup_58_payload};
  assign mulResGroup_59_valid = (inputAll_59_fork_io_outputs_0_valid && inputAll_68_fork_io_outputs_0_valid);
  assign mulResGroup_59_payload = {{7{_zz_mulResGroup_59_payload[14]}}, _zz_mulResGroup_59_payload};
  assign mulResGroup_60_valid = (inputAll_60_fork_io_outputs_0_valid && inputAll_67_fork_io_outputs_0_valid);
  assign mulResGroup_60_payload = {{6{_zz_mulResGroup_60_payload[15]}}, _zz_mulResGroup_60_payload};
  assign mulResGroup_61_valid = (inputAll_61_fork_io_outputs_0_valid && inputAll_66_fork_io_outputs_0_valid);
  assign mulResGroup_61_payload = {{6{_zz_mulResGroup_61_payload[15]}}, _zz_mulResGroup_61_payload};
  assign mulResGroup_62_valid = (inputAll_62_fork_io_outputs_0_valid && inputAll_65_fork_io_outputs_0_valid);
  assign mulResGroup_62_payload = {{5{_zz_mulResGroup_62_payload[16]}}, _zz_mulResGroup_62_payload};
  assign mulResGroup_63_valid = (inputAll_63_fork_io_outputs_0_valid && inputAll_64_fork_io_outputs_0_valid);
  assign mulResGroup_63_payload = {{5{_zz_mulResGroup_63_payload[16]}}, _zz_mulResGroup_63_payload};
  assign mulResVec_valid = ((((((((((((((((_zz_mulResVec_valid && mulResGroup_48_valid) && mulResGroup_49_valid) && mulResGroup_50_valid) && mulResGroup_51_valid) && mulResGroup_52_valid) && mulResGroup_53_valid) && mulResGroup_54_valid) && mulResGroup_55_valid) && mulResGroup_56_valid) && mulResGroup_57_valid) && mulResGroup_58_valid) && mulResGroup_59_valid) && mulResGroup_60_valid) && mulResGroup_61_valid) && mulResGroup_62_valid) && mulResGroup_63_valid);
  assign mulResGroup_0_ready = mulResVec_ready;
  assign mulResGroup_1_ready = mulResVec_ready;
  assign mulResGroup_2_ready = mulResVec_ready;
  assign mulResGroup_3_ready = mulResVec_ready;
  assign mulResGroup_4_ready = mulResVec_ready;
  assign mulResGroup_5_ready = mulResVec_ready;
  assign mulResGroup_6_ready = mulResVec_ready;
  assign mulResGroup_7_ready = mulResVec_ready;
  assign mulResGroup_8_ready = mulResVec_ready;
  assign mulResGroup_9_ready = mulResVec_ready;
  assign mulResGroup_10_ready = mulResVec_ready;
  assign mulResGroup_11_ready = mulResVec_ready;
  assign mulResGroup_12_ready = mulResVec_ready;
  assign mulResGroup_13_ready = mulResVec_ready;
  assign mulResGroup_14_ready = mulResVec_ready;
  assign mulResGroup_15_ready = mulResVec_ready;
  assign mulResGroup_16_ready = mulResVec_ready;
  assign mulResGroup_17_ready = mulResVec_ready;
  assign mulResGroup_18_ready = mulResVec_ready;
  assign mulResGroup_19_ready = mulResVec_ready;
  assign mulResGroup_20_ready = mulResVec_ready;
  assign mulResGroup_21_ready = mulResVec_ready;
  assign mulResGroup_22_ready = mulResVec_ready;
  assign mulResGroup_23_ready = mulResVec_ready;
  assign mulResGroup_24_ready = mulResVec_ready;
  assign mulResGroup_25_ready = mulResVec_ready;
  assign mulResGroup_26_ready = mulResVec_ready;
  assign mulResGroup_27_ready = mulResVec_ready;
  assign mulResGroup_28_ready = mulResVec_ready;
  assign mulResGroup_29_ready = mulResVec_ready;
  assign mulResGroup_30_ready = mulResVec_ready;
  assign mulResGroup_31_ready = mulResVec_ready;
  assign mulResGroup_32_ready = mulResVec_ready;
  assign mulResGroup_33_ready = mulResVec_ready;
  assign mulResGroup_34_ready = mulResVec_ready;
  assign mulResGroup_35_ready = mulResVec_ready;
  assign mulResGroup_36_ready = mulResVec_ready;
  assign mulResGroup_37_ready = mulResVec_ready;
  assign mulResGroup_38_ready = mulResVec_ready;
  assign mulResGroup_39_ready = mulResVec_ready;
  assign mulResGroup_40_ready = mulResVec_ready;
  assign mulResGroup_41_ready = mulResVec_ready;
  assign mulResGroup_42_ready = mulResVec_ready;
  assign mulResGroup_43_ready = mulResVec_ready;
  assign mulResGroup_44_ready = mulResVec_ready;
  assign mulResGroup_45_ready = mulResVec_ready;
  assign mulResGroup_46_ready = mulResVec_ready;
  assign mulResGroup_47_ready = mulResVec_ready;
  assign mulResGroup_48_ready = mulResVec_ready;
  assign mulResGroup_49_ready = mulResVec_ready;
  assign mulResGroup_50_ready = mulResVec_ready;
  assign mulResGroup_51_ready = mulResVec_ready;
  assign mulResGroup_52_ready = mulResVec_ready;
  assign mulResGroup_53_ready = mulResVec_ready;
  assign mulResGroup_54_ready = mulResVec_ready;
  assign mulResGroup_55_ready = mulResVec_ready;
  assign mulResGroup_56_ready = mulResVec_ready;
  assign mulResGroup_57_ready = mulResVec_ready;
  assign mulResGroup_58_ready = mulResVec_ready;
  assign mulResGroup_59_ready = mulResVec_ready;
  assign mulResGroup_60_ready = mulResVec_ready;
  assign mulResGroup_61_ready = mulResVec_ready;
  assign mulResGroup_62_ready = mulResVec_ready;
  assign mulResGroup_63_ready = mulResVec_ready;
  assign mulResVec_payload_0 = mulResGroup_0_payload;
  assign mulResVec_payload_1 = mulResGroup_1_payload;
  assign mulResVec_payload_2 = mulResGroup_2_payload;
  assign mulResVec_payload_3 = mulResGroup_3_payload;
  assign mulResVec_payload_4 = mulResGroup_4_payload;
  assign mulResVec_payload_5 = mulResGroup_5_payload;
  assign mulResVec_payload_6 = mulResGroup_6_payload;
  assign mulResVec_payload_7 = mulResGroup_7_payload;
  assign mulResVec_payload_8 = mulResGroup_8_payload;
  assign mulResVec_payload_9 = mulResGroup_9_payload;
  assign mulResVec_payload_10 = mulResGroup_10_payload;
  assign mulResVec_payload_11 = mulResGroup_11_payload;
  assign mulResVec_payload_12 = mulResGroup_12_payload;
  assign mulResVec_payload_13 = mulResGroup_13_payload;
  assign mulResVec_payload_14 = mulResGroup_14_payload;
  assign mulResVec_payload_15 = mulResGroup_15_payload;
  assign mulResVec_payload_16 = mulResGroup_16_payload;
  assign mulResVec_payload_17 = mulResGroup_17_payload;
  assign mulResVec_payload_18 = mulResGroup_18_payload;
  assign mulResVec_payload_19 = mulResGroup_19_payload;
  assign mulResVec_payload_20 = mulResGroup_20_payload;
  assign mulResVec_payload_21 = mulResGroup_21_payload;
  assign mulResVec_payload_22 = mulResGroup_22_payload;
  assign mulResVec_payload_23 = mulResGroup_23_payload;
  assign mulResVec_payload_24 = mulResGroup_24_payload;
  assign mulResVec_payload_25 = mulResGroup_25_payload;
  assign mulResVec_payload_26 = mulResGroup_26_payload;
  assign mulResVec_payload_27 = mulResGroup_27_payload;
  assign mulResVec_payload_28 = mulResGroup_28_payload;
  assign mulResVec_payload_29 = mulResGroup_29_payload;
  assign mulResVec_payload_30 = mulResGroup_30_payload;
  assign mulResVec_payload_31 = mulResGroup_31_payload;
  assign mulResVec_payload_32 = mulResGroup_32_payload;
  assign mulResVec_payload_33 = mulResGroup_33_payload;
  assign mulResVec_payload_34 = mulResGroup_34_payload;
  assign mulResVec_payload_35 = mulResGroup_35_payload;
  assign mulResVec_payload_36 = mulResGroup_36_payload;
  assign mulResVec_payload_37 = mulResGroup_37_payload;
  assign mulResVec_payload_38 = mulResGroup_38_payload;
  assign mulResVec_payload_39 = mulResGroup_39_payload;
  assign mulResVec_payload_40 = mulResGroup_40_payload;
  assign mulResVec_payload_41 = mulResGroup_41_payload;
  assign mulResVec_payload_42 = mulResGroup_42_payload;
  assign mulResVec_payload_43 = mulResGroup_43_payload;
  assign mulResVec_payload_44 = mulResGroup_44_payload;
  assign mulResVec_payload_45 = mulResGroup_45_payload;
  assign mulResVec_payload_46 = mulResGroup_46_payload;
  assign mulResVec_payload_47 = mulResGroup_47_payload;
  assign mulResVec_payload_48 = mulResGroup_48_payload;
  assign mulResVec_payload_49 = mulResGroup_49_payload;
  assign mulResVec_payload_50 = mulResGroup_50_payload;
  assign mulResVec_payload_51 = mulResGroup_51_payload;
  assign mulResVec_payload_52 = mulResGroup_52_payload;
  assign mulResVec_payload_53 = mulResGroup_53_payload;
  assign mulResVec_payload_54 = mulResGroup_54_payload;
  assign mulResVec_payload_55 = mulResGroup_55_payload;
  assign mulResVec_payload_56 = mulResGroup_56_payload;
  assign mulResVec_payload_57 = mulResGroup_57_payload;
  assign mulResVec_payload_58 = mulResGroup_58_payload;
  assign mulResVec_payload_59 = mulResGroup_59_payload;
  assign mulResVec_payload_60 = mulResGroup_60_payload;
  assign mulResVec_payload_61 = mulResGroup_61_payload;
  assign mulResVec_payload_62 = mulResGroup_62_payload;
  assign mulResVec_payload_63 = mulResGroup_63_payload;
  assign mulResVec_translated_valid = mulResVec_valid;
  assign mulResVec_ready = mulResVec_translated_ready;
  assign mulResVec_translated_payload = ($signed(_zz_mulResVec_translated_payload) + $signed(_zz_mulResVec_translated_payload_31));
  assign io_output_valid = mulResVec_translated_valid;
  assign mulResVec_translated_ready = io_output_ready;
  assign io_output_payload = mulResVec_translated_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      inputAll_0_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_1_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_2_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_3_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_4_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_5_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_6_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_7_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_8_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_9_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_10_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_11_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_12_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_13_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_14_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_15_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_16_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_17_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_18_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_19_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_20_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_21_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_22_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_23_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_24_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_25_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_26_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_27_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_28_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_29_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_30_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_31_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_32_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_33_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_34_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_35_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_36_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_37_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_38_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_39_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_40_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_41_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_42_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_43_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_44_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_45_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_46_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_47_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_48_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_49_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_50_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_51_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_52_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_53_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_54_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_55_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_56_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_57_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_58_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_59_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_60_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_61_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_62_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_63_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_64_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_65_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_66_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_67_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_68_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_69_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_70_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_71_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_72_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_73_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_74_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_75_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_76_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_77_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_78_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_79_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_80_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_81_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_82_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_83_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_84_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_85_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_86_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_87_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_88_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_89_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_90_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_91_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_92_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_93_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_94_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_95_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_96_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_97_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_98_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_99_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_100_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_101_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_102_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_103_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_104_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_105_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_106_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_107_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_108_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_109_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_110_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_111_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_112_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_113_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_114_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_115_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_116_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_117_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_118_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_119_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_120_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_121_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_122_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_123_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_124_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_125_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_126_fork_io_outputs_1_rValid <= 1'b0;
      inputAll_127_fork_io_outputs_1_rValid <= 1'b0;
    end else begin
      if(inputAll_0_fork_io_outputs_1_ready) begin
        inputAll_0_fork_io_outputs_1_rValid <= inputAll_0_fork_io_outputs_1_valid;
      end
      if(inputAll_1_fork_io_outputs_1_ready) begin
        inputAll_1_fork_io_outputs_1_rValid <= inputAll_1_fork_io_outputs_1_valid;
      end
      if(inputAll_2_fork_io_outputs_1_ready) begin
        inputAll_2_fork_io_outputs_1_rValid <= inputAll_2_fork_io_outputs_1_valid;
      end
      if(inputAll_3_fork_io_outputs_1_ready) begin
        inputAll_3_fork_io_outputs_1_rValid <= inputAll_3_fork_io_outputs_1_valid;
      end
      if(inputAll_4_fork_io_outputs_1_ready) begin
        inputAll_4_fork_io_outputs_1_rValid <= inputAll_4_fork_io_outputs_1_valid;
      end
      if(inputAll_5_fork_io_outputs_1_ready) begin
        inputAll_5_fork_io_outputs_1_rValid <= inputAll_5_fork_io_outputs_1_valid;
      end
      if(inputAll_6_fork_io_outputs_1_ready) begin
        inputAll_6_fork_io_outputs_1_rValid <= inputAll_6_fork_io_outputs_1_valid;
      end
      if(inputAll_7_fork_io_outputs_1_ready) begin
        inputAll_7_fork_io_outputs_1_rValid <= inputAll_7_fork_io_outputs_1_valid;
      end
      if(inputAll_8_fork_io_outputs_1_ready) begin
        inputAll_8_fork_io_outputs_1_rValid <= inputAll_8_fork_io_outputs_1_valid;
      end
      if(inputAll_9_fork_io_outputs_1_ready) begin
        inputAll_9_fork_io_outputs_1_rValid <= inputAll_9_fork_io_outputs_1_valid;
      end
      if(inputAll_10_fork_io_outputs_1_ready) begin
        inputAll_10_fork_io_outputs_1_rValid <= inputAll_10_fork_io_outputs_1_valid;
      end
      if(inputAll_11_fork_io_outputs_1_ready) begin
        inputAll_11_fork_io_outputs_1_rValid <= inputAll_11_fork_io_outputs_1_valid;
      end
      if(inputAll_12_fork_io_outputs_1_ready) begin
        inputAll_12_fork_io_outputs_1_rValid <= inputAll_12_fork_io_outputs_1_valid;
      end
      if(inputAll_13_fork_io_outputs_1_ready) begin
        inputAll_13_fork_io_outputs_1_rValid <= inputAll_13_fork_io_outputs_1_valid;
      end
      if(inputAll_14_fork_io_outputs_1_ready) begin
        inputAll_14_fork_io_outputs_1_rValid <= inputAll_14_fork_io_outputs_1_valid;
      end
      if(inputAll_15_fork_io_outputs_1_ready) begin
        inputAll_15_fork_io_outputs_1_rValid <= inputAll_15_fork_io_outputs_1_valid;
      end
      if(inputAll_16_fork_io_outputs_1_ready) begin
        inputAll_16_fork_io_outputs_1_rValid <= inputAll_16_fork_io_outputs_1_valid;
      end
      if(inputAll_17_fork_io_outputs_1_ready) begin
        inputAll_17_fork_io_outputs_1_rValid <= inputAll_17_fork_io_outputs_1_valid;
      end
      if(inputAll_18_fork_io_outputs_1_ready) begin
        inputAll_18_fork_io_outputs_1_rValid <= inputAll_18_fork_io_outputs_1_valid;
      end
      if(inputAll_19_fork_io_outputs_1_ready) begin
        inputAll_19_fork_io_outputs_1_rValid <= inputAll_19_fork_io_outputs_1_valid;
      end
      if(inputAll_20_fork_io_outputs_1_ready) begin
        inputAll_20_fork_io_outputs_1_rValid <= inputAll_20_fork_io_outputs_1_valid;
      end
      if(inputAll_21_fork_io_outputs_1_ready) begin
        inputAll_21_fork_io_outputs_1_rValid <= inputAll_21_fork_io_outputs_1_valid;
      end
      if(inputAll_22_fork_io_outputs_1_ready) begin
        inputAll_22_fork_io_outputs_1_rValid <= inputAll_22_fork_io_outputs_1_valid;
      end
      if(inputAll_23_fork_io_outputs_1_ready) begin
        inputAll_23_fork_io_outputs_1_rValid <= inputAll_23_fork_io_outputs_1_valid;
      end
      if(inputAll_24_fork_io_outputs_1_ready) begin
        inputAll_24_fork_io_outputs_1_rValid <= inputAll_24_fork_io_outputs_1_valid;
      end
      if(inputAll_25_fork_io_outputs_1_ready) begin
        inputAll_25_fork_io_outputs_1_rValid <= inputAll_25_fork_io_outputs_1_valid;
      end
      if(inputAll_26_fork_io_outputs_1_ready) begin
        inputAll_26_fork_io_outputs_1_rValid <= inputAll_26_fork_io_outputs_1_valid;
      end
      if(inputAll_27_fork_io_outputs_1_ready) begin
        inputAll_27_fork_io_outputs_1_rValid <= inputAll_27_fork_io_outputs_1_valid;
      end
      if(inputAll_28_fork_io_outputs_1_ready) begin
        inputAll_28_fork_io_outputs_1_rValid <= inputAll_28_fork_io_outputs_1_valid;
      end
      if(inputAll_29_fork_io_outputs_1_ready) begin
        inputAll_29_fork_io_outputs_1_rValid <= inputAll_29_fork_io_outputs_1_valid;
      end
      if(inputAll_30_fork_io_outputs_1_ready) begin
        inputAll_30_fork_io_outputs_1_rValid <= inputAll_30_fork_io_outputs_1_valid;
      end
      if(inputAll_31_fork_io_outputs_1_ready) begin
        inputAll_31_fork_io_outputs_1_rValid <= inputAll_31_fork_io_outputs_1_valid;
      end
      if(inputAll_32_fork_io_outputs_1_ready) begin
        inputAll_32_fork_io_outputs_1_rValid <= inputAll_32_fork_io_outputs_1_valid;
      end
      if(inputAll_33_fork_io_outputs_1_ready) begin
        inputAll_33_fork_io_outputs_1_rValid <= inputAll_33_fork_io_outputs_1_valid;
      end
      if(inputAll_34_fork_io_outputs_1_ready) begin
        inputAll_34_fork_io_outputs_1_rValid <= inputAll_34_fork_io_outputs_1_valid;
      end
      if(inputAll_35_fork_io_outputs_1_ready) begin
        inputAll_35_fork_io_outputs_1_rValid <= inputAll_35_fork_io_outputs_1_valid;
      end
      if(inputAll_36_fork_io_outputs_1_ready) begin
        inputAll_36_fork_io_outputs_1_rValid <= inputAll_36_fork_io_outputs_1_valid;
      end
      if(inputAll_37_fork_io_outputs_1_ready) begin
        inputAll_37_fork_io_outputs_1_rValid <= inputAll_37_fork_io_outputs_1_valid;
      end
      if(inputAll_38_fork_io_outputs_1_ready) begin
        inputAll_38_fork_io_outputs_1_rValid <= inputAll_38_fork_io_outputs_1_valid;
      end
      if(inputAll_39_fork_io_outputs_1_ready) begin
        inputAll_39_fork_io_outputs_1_rValid <= inputAll_39_fork_io_outputs_1_valid;
      end
      if(inputAll_40_fork_io_outputs_1_ready) begin
        inputAll_40_fork_io_outputs_1_rValid <= inputAll_40_fork_io_outputs_1_valid;
      end
      if(inputAll_41_fork_io_outputs_1_ready) begin
        inputAll_41_fork_io_outputs_1_rValid <= inputAll_41_fork_io_outputs_1_valid;
      end
      if(inputAll_42_fork_io_outputs_1_ready) begin
        inputAll_42_fork_io_outputs_1_rValid <= inputAll_42_fork_io_outputs_1_valid;
      end
      if(inputAll_43_fork_io_outputs_1_ready) begin
        inputAll_43_fork_io_outputs_1_rValid <= inputAll_43_fork_io_outputs_1_valid;
      end
      if(inputAll_44_fork_io_outputs_1_ready) begin
        inputAll_44_fork_io_outputs_1_rValid <= inputAll_44_fork_io_outputs_1_valid;
      end
      if(inputAll_45_fork_io_outputs_1_ready) begin
        inputAll_45_fork_io_outputs_1_rValid <= inputAll_45_fork_io_outputs_1_valid;
      end
      if(inputAll_46_fork_io_outputs_1_ready) begin
        inputAll_46_fork_io_outputs_1_rValid <= inputAll_46_fork_io_outputs_1_valid;
      end
      if(inputAll_47_fork_io_outputs_1_ready) begin
        inputAll_47_fork_io_outputs_1_rValid <= inputAll_47_fork_io_outputs_1_valid;
      end
      if(inputAll_48_fork_io_outputs_1_ready) begin
        inputAll_48_fork_io_outputs_1_rValid <= inputAll_48_fork_io_outputs_1_valid;
      end
      if(inputAll_49_fork_io_outputs_1_ready) begin
        inputAll_49_fork_io_outputs_1_rValid <= inputAll_49_fork_io_outputs_1_valid;
      end
      if(inputAll_50_fork_io_outputs_1_ready) begin
        inputAll_50_fork_io_outputs_1_rValid <= inputAll_50_fork_io_outputs_1_valid;
      end
      if(inputAll_51_fork_io_outputs_1_ready) begin
        inputAll_51_fork_io_outputs_1_rValid <= inputAll_51_fork_io_outputs_1_valid;
      end
      if(inputAll_52_fork_io_outputs_1_ready) begin
        inputAll_52_fork_io_outputs_1_rValid <= inputAll_52_fork_io_outputs_1_valid;
      end
      if(inputAll_53_fork_io_outputs_1_ready) begin
        inputAll_53_fork_io_outputs_1_rValid <= inputAll_53_fork_io_outputs_1_valid;
      end
      if(inputAll_54_fork_io_outputs_1_ready) begin
        inputAll_54_fork_io_outputs_1_rValid <= inputAll_54_fork_io_outputs_1_valid;
      end
      if(inputAll_55_fork_io_outputs_1_ready) begin
        inputAll_55_fork_io_outputs_1_rValid <= inputAll_55_fork_io_outputs_1_valid;
      end
      if(inputAll_56_fork_io_outputs_1_ready) begin
        inputAll_56_fork_io_outputs_1_rValid <= inputAll_56_fork_io_outputs_1_valid;
      end
      if(inputAll_57_fork_io_outputs_1_ready) begin
        inputAll_57_fork_io_outputs_1_rValid <= inputAll_57_fork_io_outputs_1_valid;
      end
      if(inputAll_58_fork_io_outputs_1_ready) begin
        inputAll_58_fork_io_outputs_1_rValid <= inputAll_58_fork_io_outputs_1_valid;
      end
      if(inputAll_59_fork_io_outputs_1_ready) begin
        inputAll_59_fork_io_outputs_1_rValid <= inputAll_59_fork_io_outputs_1_valid;
      end
      if(inputAll_60_fork_io_outputs_1_ready) begin
        inputAll_60_fork_io_outputs_1_rValid <= inputAll_60_fork_io_outputs_1_valid;
      end
      if(inputAll_61_fork_io_outputs_1_ready) begin
        inputAll_61_fork_io_outputs_1_rValid <= inputAll_61_fork_io_outputs_1_valid;
      end
      if(inputAll_62_fork_io_outputs_1_ready) begin
        inputAll_62_fork_io_outputs_1_rValid <= inputAll_62_fork_io_outputs_1_valid;
      end
      if(inputAll_63_fork_io_outputs_1_ready) begin
        inputAll_63_fork_io_outputs_1_rValid <= inputAll_63_fork_io_outputs_1_valid;
      end
      if(inputAll_64_fork_io_outputs_1_ready) begin
        inputAll_64_fork_io_outputs_1_rValid <= inputAll_64_fork_io_outputs_1_valid;
      end
      if(inputAll_65_fork_io_outputs_1_ready) begin
        inputAll_65_fork_io_outputs_1_rValid <= inputAll_65_fork_io_outputs_1_valid;
      end
      if(inputAll_66_fork_io_outputs_1_ready) begin
        inputAll_66_fork_io_outputs_1_rValid <= inputAll_66_fork_io_outputs_1_valid;
      end
      if(inputAll_67_fork_io_outputs_1_ready) begin
        inputAll_67_fork_io_outputs_1_rValid <= inputAll_67_fork_io_outputs_1_valid;
      end
      if(inputAll_68_fork_io_outputs_1_ready) begin
        inputAll_68_fork_io_outputs_1_rValid <= inputAll_68_fork_io_outputs_1_valid;
      end
      if(inputAll_69_fork_io_outputs_1_ready) begin
        inputAll_69_fork_io_outputs_1_rValid <= inputAll_69_fork_io_outputs_1_valid;
      end
      if(inputAll_70_fork_io_outputs_1_ready) begin
        inputAll_70_fork_io_outputs_1_rValid <= inputAll_70_fork_io_outputs_1_valid;
      end
      if(inputAll_71_fork_io_outputs_1_ready) begin
        inputAll_71_fork_io_outputs_1_rValid <= inputAll_71_fork_io_outputs_1_valid;
      end
      if(inputAll_72_fork_io_outputs_1_ready) begin
        inputAll_72_fork_io_outputs_1_rValid <= inputAll_72_fork_io_outputs_1_valid;
      end
      if(inputAll_73_fork_io_outputs_1_ready) begin
        inputAll_73_fork_io_outputs_1_rValid <= inputAll_73_fork_io_outputs_1_valid;
      end
      if(inputAll_74_fork_io_outputs_1_ready) begin
        inputAll_74_fork_io_outputs_1_rValid <= inputAll_74_fork_io_outputs_1_valid;
      end
      if(inputAll_75_fork_io_outputs_1_ready) begin
        inputAll_75_fork_io_outputs_1_rValid <= inputAll_75_fork_io_outputs_1_valid;
      end
      if(inputAll_76_fork_io_outputs_1_ready) begin
        inputAll_76_fork_io_outputs_1_rValid <= inputAll_76_fork_io_outputs_1_valid;
      end
      if(inputAll_77_fork_io_outputs_1_ready) begin
        inputAll_77_fork_io_outputs_1_rValid <= inputAll_77_fork_io_outputs_1_valid;
      end
      if(inputAll_78_fork_io_outputs_1_ready) begin
        inputAll_78_fork_io_outputs_1_rValid <= inputAll_78_fork_io_outputs_1_valid;
      end
      if(inputAll_79_fork_io_outputs_1_ready) begin
        inputAll_79_fork_io_outputs_1_rValid <= inputAll_79_fork_io_outputs_1_valid;
      end
      if(inputAll_80_fork_io_outputs_1_ready) begin
        inputAll_80_fork_io_outputs_1_rValid <= inputAll_80_fork_io_outputs_1_valid;
      end
      if(inputAll_81_fork_io_outputs_1_ready) begin
        inputAll_81_fork_io_outputs_1_rValid <= inputAll_81_fork_io_outputs_1_valid;
      end
      if(inputAll_82_fork_io_outputs_1_ready) begin
        inputAll_82_fork_io_outputs_1_rValid <= inputAll_82_fork_io_outputs_1_valid;
      end
      if(inputAll_83_fork_io_outputs_1_ready) begin
        inputAll_83_fork_io_outputs_1_rValid <= inputAll_83_fork_io_outputs_1_valid;
      end
      if(inputAll_84_fork_io_outputs_1_ready) begin
        inputAll_84_fork_io_outputs_1_rValid <= inputAll_84_fork_io_outputs_1_valid;
      end
      if(inputAll_85_fork_io_outputs_1_ready) begin
        inputAll_85_fork_io_outputs_1_rValid <= inputAll_85_fork_io_outputs_1_valid;
      end
      if(inputAll_86_fork_io_outputs_1_ready) begin
        inputAll_86_fork_io_outputs_1_rValid <= inputAll_86_fork_io_outputs_1_valid;
      end
      if(inputAll_87_fork_io_outputs_1_ready) begin
        inputAll_87_fork_io_outputs_1_rValid <= inputAll_87_fork_io_outputs_1_valid;
      end
      if(inputAll_88_fork_io_outputs_1_ready) begin
        inputAll_88_fork_io_outputs_1_rValid <= inputAll_88_fork_io_outputs_1_valid;
      end
      if(inputAll_89_fork_io_outputs_1_ready) begin
        inputAll_89_fork_io_outputs_1_rValid <= inputAll_89_fork_io_outputs_1_valid;
      end
      if(inputAll_90_fork_io_outputs_1_ready) begin
        inputAll_90_fork_io_outputs_1_rValid <= inputAll_90_fork_io_outputs_1_valid;
      end
      if(inputAll_91_fork_io_outputs_1_ready) begin
        inputAll_91_fork_io_outputs_1_rValid <= inputAll_91_fork_io_outputs_1_valid;
      end
      if(inputAll_92_fork_io_outputs_1_ready) begin
        inputAll_92_fork_io_outputs_1_rValid <= inputAll_92_fork_io_outputs_1_valid;
      end
      if(inputAll_93_fork_io_outputs_1_ready) begin
        inputAll_93_fork_io_outputs_1_rValid <= inputAll_93_fork_io_outputs_1_valid;
      end
      if(inputAll_94_fork_io_outputs_1_ready) begin
        inputAll_94_fork_io_outputs_1_rValid <= inputAll_94_fork_io_outputs_1_valid;
      end
      if(inputAll_95_fork_io_outputs_1_ready) begin
        inputAll_95_fork_io_outputs_1_rValid <= inputAll_95_fork_io_outputs_1_valid;
      end
      if(inputAll_96_fork_io_outputs_1_ready) begin
        inputAll_96_fork_io_outputs_1_rValid <= inputAll_96_fork_io_outputs_1_valid;
      end
      if(inputAll_97_fork_io_outputs_1_ready) begin
        inputAll_97_fork_io_outputs_1_rValid <= inputAll_97_fork_io_outputs_1_valid;
      end
      if(inputAll_98_fork_io_outputs_1_ready) begin
        inputAll_98_fork_io_outputs_1_rValid <= inputAll_98_fork_io_outputs_1_valid;
      end
      if(inputAll_99_fork_io_outputs_1_ready) begin
        inputAll_99_fork_io_outputs_1_rValid <= inputAll_99_fork_io_outputs_1_valid;
      end
      if(inputAll_100_fork_io_outputs_1_ready) begin
        inputAll_100_fork_io_outputs_1_rValid <= inputAll_100_fork_io_outputs_1_valid;
      end
      if(inputAll_101_fork_io_outputs_1_ready) begin
        inputAll_101_fork_io_outputs_1_rValid <= inputAll_101_fork_io_outputs_1_valid;
      end
      if(inputAll_102_fork_io_outputs_1_ready) begin
        inputAll_102_fork_io_outputs_1_rValid <= inputAll_102_fork_io_outputs_1_valid;
      end
      if(inputAll_103_fork_io_outputs_1_ready) begin
        inputAll_103_fork_io_outputs_1_rValid <= inputAll_103_fork_io_outputs_1_valid;
      end
      if(inputAll_104_fork_io_outputs_1_ready) begin
        inputAll_104_fork_io_outputs_1_rValid <= inputAll_104_fork_io_outputs_1_valid;
      end
      if(inputAll_105_fork_io_outputs_1_ready) begin
        inputAll_105_fork_io_outputs_1_rValid <= inputAll_105_fork_io_outputs_1_valid;
      end
      if(inputAll_106_fork_io_outputs_1_ready) begin
        inputAll_106_fork_io_outputs_1_rValid <= inputAll_106_fork_io_outputs_1_valid;
      end
      if(inputAll_107_fork_io_outputs_1_ready) begin
        inputAll_107_fork_io_outputs_1_rValid <= inputAll_107_fork_io_outputs_1_valid;
      end
      if(inputAll_108_fork_io_outputs_1_ready) begin
        inputAll_108_fork_io_outputs_1_rValid <= inputAll_108_fork_io_outputs_1_valid;
      end
      if(inputAll_109_fork_io_outputs_1_ready) begin
        inputAll_109_fork_io_outputs_1_rValid <= inputAll_109_fork_io_outputs_1_valid;
      end
      if(inputAll_110_fork_io_outputs_1_ready) begin
        inputAll_110_fork_io_outputs_1_rValid <= inputAll_110_fork_io_outputs_1_valid;
      end
      if(inputAll_111_fork_io_outputs_1_ready) begin
        inputAll_111_fork_io_outputs_1_rValid <= inputAll_111_fork_io_outputs_1_valid;
      end
      if(inputAll_112_fork_io_outputs_1_ready) begin
        inputAll_112_fork_io_outputs_1_rValid <= inputAll_112_fork_io_outputs_1_valid;
      end
      if(inputAll_113_fork_io_outputs_1_ready) begin
        inputAll_113_fork_io_outputs_1_rValid <= inputAll_113_fork_io_outputs_1_valid;
      end
      if(inputAll_114_fork_io_outputs_1_ready) begin
        inputAll_114_fork_io_outputs_1_rValid <= inputAll_114_fork_io_outputs_1_valid;
      end
      if(inputAll_115_fork_io_outputs_1_ready) begin
        inputAll_115_fork_io_outputs_1_rValid <= inputAll_115_fork_io_outputs_1_valid;
      end
      if(inputAll_116_fork_io_outputs_1_ready) begin
        inputAll_116_fork_io_outputs_1_rValid <= inputAll_116_fork_io_outputs_1_valid;
      end
      if(inputAll_117_fork_io_outputs_1_ready) begin
        inputAll_117_fork_io_outputs_1_rValid <= inputAll_117_fork_io_outputs_1_valid;
      end
      if(inputAll_118_fork_io_outputs_1_ready) begin
        inputAll_118_fork_io_outputs_1_rValid <= inputAll_118_fork_io_outputs_1_valid;
      end
      if(inputAll_119_fork_io_outputs_1_ready) begin
        inputAll_119_fork_io_outputs_1_rValid <= inputAll_119_fork_io_outputs_1_valid;
      end
      if(inputAll_120_fork_io_outputs_1_ready) begin
        inputAll_120_fork_io_outputs_1_rValid <= inputAll_120_fork_io_outputs_1_valid;
      end
      if(inputAll_121_fork_io_outputs_1_ready) begin
        inputAll_121_fork_io_outputs_1_rValid <= inputAll_121_fork_io_outputs_1_valid;
      end
      if(inputAll_122_fork_io_outputs_1_ready) begin
        inputAll_122_fork_io_outputs_1_rValid <= inputAll_122_fork_io_outputs_1_valid;
      end
      if(inputAll_123_fork_io_outputs_1_ready) begin
        inputAll_123_fork_io_outputs_1_rValid <= inputAll_123_fork_io_outputs_1_valid;
      end
      if(inputAll_124_fork_io_outputs_1_ready) begin
        inputAll_124_fork_io_outputs_1_rValid <= inputAll_124_fork_io_outputs_1_valid;
      end
      if(inputAll_125_fork_io_outputs_1_ready) begin
        inputAll_125_fork_io_outputs_1_rValid <= inputAll_125_fork_io_outputs_1_valid;
      end
      if(inputAll_126_fork_io_outputs_1_ready) begin
        inputAll_126_fork_io_outputs_1_rValid <= inputAll_126_fork_io_outputs_1_valid;
      end
      if(inputAll_127_fork_io_outputs_1_ready) begin
        inputAll_127_fork_io_outputs_1_rValid <= inputAll_127_fork_io_outputs_1_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(inputAll_0_fork_io_outputs_1_ready) begin
      inputAll_0_fork_io_outputs_1_rData <= inputAll_0_fork_io_outputs_1_payload;
    end
    if(inputAll_1_fork_io_outputs_1_ready) begin
      inputAll_1_fork_io_outputs_1_rData <= inputAll_1_fork_io_outputs_1_payload;
    end
    if(inputAll_2_fork_io_outputs_1_ready) begin
      inputAll_2_fork_io_outputs_1_rData <= inputAll_2_fork_io_outputs_1_payload;
    end
    if(inputAll_3_fork_io_outputs_1_ready) begin
      inputAll_3_fork_io_outputs_1_rData <= inputAll_3_fork_io_outputs_1_payload;
    end
    if(inputAll_4_fork_io_outputs_1_ready) begin
      inputAll_4_fork_io_outputs_1_rData <= inputAll_4_fork_io_outputs_1_payload;
    end
    if(inputAll_5_fork_io_outputs_1_ready) begin
      inputAll_5_fork_io_outputs_1_rData <= inputAll_5_fork_io_outputs_1_payload;
    end
    if(inputAll_6_fork_io_outputs_1_ready) begin
      inputAll_6_fork_io_outputs_1_rData <= inputAll_6_fork_io_outputs_1_payload;
    end
    if(inputAll_7_fork_io_outputs_1_ready) begin
      inputAll_7_fork_io_outputs_1_rData <= inputAll_7_fork_io_outputs_1_payload;
    end
    if(inputAll_8_fork_io_outputs_1_ready) begin
      inputAll_8_fork_io_outputs_1_rData <= inputAll_8_fork_io_outputs_1_payload;
    end
    if(inputAll_9_fork_io_outputs_1_ready) begin
      inputAll_9_fork_io_outputs_1_rData <= inputAll_9_fork_io_outputs_1_payload;
    end
    if(inputAll_10_fork_io_outputs_1_ready) begin
      inputAll_10_fork_io_outputs_1_rData <= inputAll_10_fork_io_outputs_1_payload;
    end
    if(inputAll_11_fork_io_outputs_1_ready) begin
      inputAll_11_fork_io_outputs_1_rData <= inputAll_11_fork_io_outputs_1_payload;
    end
    if(inputAll_12_fork_io_outputs_1_ready) begin
      inputAll_12_fork_io_outputs_1_rData <= inputAll_12_fork_io_outputs_1_payload;
    end
    if(inputAll_13_fork_io_outputs_1_ready) begin
      inputAll_13_fork_io_outputs_1_rData <= inputAll_13_fork_io_outputs_1_payload;
    end
    if(inputAll_14_fork_io_outputs_1_ready) begin
      inputAll_14_fork_io_outputs_1_rData <= inputAll_14_fork_io_outputs_1_payload;
    end
    if(inputAll_15_fork_io_outputs_1_ready) begin
      inputAll_15_fork_io_outputs_1_rData <= inputAll_15_fork_io_outputs_1_payload;
    end
    if(inputAll_16_fork_io_outputs_1_ready) begin
      inputAll_16_fork_io_outputs_1_rData <= inputAll_16_fork_io_outputs_1_payload;
    end
    if(inputAll_17_fork_io_outputs_1_ready) begin
      inputAll_17_fork_io_outputs_1_rData <= inputAll_17_fork_io_outputs_1_payload;
    end
    if(inputAll_18_fork_io_outputs_1_ready) begin
      inputAll_18_fork_io_outputs_1_rData <= inputAll_18_fork_io_outputs_1_payload;
    end
    if(inputAll_19_fork_io_outputs_1_ready) begin
      inputAll_19_fork_io_outputs_1_rData <= inputAll_19_fork_io_outputs_1_payload;
    end
    if(inputAll_20_fork_io_outputs_1_ready) begin
      inputAll_20_fork_io_outputs_1_rData <= inputAll_20_fork_io_outputs_1_payload;
    end
    if(inputAll_21_fork_io_outputs_1_ready) begin
      inputAll_21_fork_io_outputs_1_rData <= inputAll_21_fork_io_outputs_1_payload;
    end
    if(inputAll_22_fork_io_outputs_1_ready) begin
      inputAll_22_fork_io_outputs_1_rData <= inputAll_22_fork_io_outputs_1_payload;
    end
    if(inputAll_23_fork_io_outputs_1_ready) begin
      inputAll_23_fork_io_outputs_1_rData <= inputAll_23_fork_io_outputs_1_payload;
    end
    if(inputAll_24_fork_io_outputs_1_ready) begin
      inputAll_24_fork_io_outputs_1_rData <= inputAll_24_fork_io_outputs_1_payload;
    end
    if(inputAll_25_fork_io_outputs_1_ready) begin
      inputAll_25_fork_io_outputs_1_rData <= inputAll_25_fork_io_outputs_1_payload;
    end
    if(inputAll_26_fork_io_outputs_1_ready) begin
      inputAll_26_fork_io_outputs_1_rData <= inputAll_26_fork_io_outputs_1_payload;
    end
    if(inputAll_27_fork_io_outputs_1_ready) begin
      inputAll_27_fork_io_outputs_1_rData <= inputAll_27_fork_io_outputs_1_payload;
    end
    if(inputAll_28_fork_io_outputs_1_ready) begin
      inputAll_28_fork_io_outputs_1_rData <= inputAll_28_fork_io_outputs_1_payload;
    end
    if(inputAll_29_fork_io_outputs_1_ready) begin
      inputAll_29_fork_io_outputs_1_rData <= inputAll_29_fork_io_outputs_1_payload;
    end
    if(inputAll_30_fork_io_outputs_1_ready) begin
      inputAll_30_fork_io_outputs_1_rData <= inputAll_30_fork_io_outputs_1_payload;
    end
    if(inputAll_31_fork_io_outputs_1_ready) begin
      inputAll_31_fork_io_outputs_1_rData <= inputAll_31_fork_io_outputs_1_payload;
    end
    if(inputAll_32_fork_io_outputs_1_ready) begin
      inputAll_32_fork_io_outputs_1_rData <= inputAll_32_fork_io_outputs_1_payload;
    end
    if(inputAll_33_fork_io_outputs_1_ready) begin
      inputAll_33_fork_io_outputs_1_rData <= inputAll_33_fork_io_outputs_1_payload;
    end
    if(inputAll_34_fork_io_outputs_1_ready) begin
      inputAll_34_fork_io_outputs_1_rData <= inputAll_34_fork_io_outputs_1_payload;
    end
    if(inputAll_35_fork_io_outputs_1_ready) begin
      inputAll_35_fork_io_outputs_1_rData <= inputAll_35_fork_io_outputs_1_payload;
    end
    if(inputAll_36_fork_io_outputs_1_ready) begin
      inputAll_36_fork_io_outputs_1_rData <= inputAll_36_fork_io_outputs_1_payload;
    end
    if(inputAll_37_fork_io_outputs_1_ready) begin
      inputAll_37_fork_io_outputs_1_rData <= inputAll_37_fork_io_outputs_1_payload;
    end
    if(inputAll_38_fork_io_outputs_1_ready) begin
      inputAll_38_fork_io_outputs_1_rData <= inputAll_38_fork_io_outputs_1_payload;
    end
    if(inputAll_39_fork_io_outputs_1_ready) begin
      inputAll_39_fork_io_outputs_1_rData <= inputAll_39_fork_io_outputs_1_payload;
    end
    if(inputAll_40_fork_io_outputs_1_ready) begin
      inputAll_40_fork_io_outputs_1_rData <= inputAll_40_fork_io_outputs_1_payload;
    end
    if(inputAll_41_fork_io_outputs_1_ready) begin
      inputAll_41_fork_io_outputs_1_rData <= inputAll_41_fork_io_outputs_1_payload;
    end
    if(inputAll_42_fork_io_outputs_1_ready) begin
      inputAll_42_fork_io_outputs_1_rData <= inputAll_42_fork_io_outputs_1_payload;
    end
    if(inputAll_43_fork_io_outputs_1_ready) begin
      inputAll_43_fork_io_outputs_1_rData <= inputAll_43_fork_io_outputs_1_payload;
    end
    if(inputAll_44_fork_io_outputs_1_ready) begin
      inputAll_44_fork_io_outputs_1_rData <= inputAll_44_fork_io_outputs_1_payload;
    end
    if(inputAll_45_fork_io_outputs_1_ready) begin
      inputAll_45_fork_io_outputs_1_rData <= inputAll_45_fork_io_outputs_1_payload;
    end
    if(inputAll_46_fork_io_outputs_1_ready) begin
      inputAll_46_fork_io_outputs_1_rData <= inputAll_46_fork_io_outputs_1_payload;
    end
    if(inputAll_47_fork_io_outputs_1_ready) begin
      inputAll_47_fork_io_outputs_1_rData <= inputAll_47_fork_io_outputs_1_payload;
    end
    if(inputAll_48_fork_io_outputs_1_ready) begin
      inputAll_48_fork_io_outputs_1_rData <= inputAll_48_fork_io_outputs_1_payload;
    end
    if(inputAll_49_fork_io_outputs_1_ready) begin
      inputAll_49_fork_io_outputs_1_rData <= inputAll_49_fork_io_outputs_1_payload;
    end
    if(inputAll_50_fork_io_outputs_1_ready) begin
      inputAll_50_fork_io_outputs_1_rData <= inputAll_50_fork_io_outputs_1_payload;
    end
    if(inputAll_51_fork_io_outputs_1_ready) begin
      inputAll_51_fork_io_outputs_1_rData <= inputAll_51_fork_io_outputs_1_payload;
    end
    if(inputAll_52_fork_io_outputs_1_ready) begin
      inputAll_52_fork_io_outputs_1_rData <= inputAll_52_fork_io_outputs_1_payload;
    end
    if(inputAll_53_fork_io_outputs_1_ready) begin
      inputAll_53_fork_io_outputs_1_rData <= inputAll_53_fork_io_outputs_1_payload;
    end
    if(inputAll_54_fork_io_outputs_1_ready) begin
      inputAll_54_fork_io_outputs_1_rData <= inputAll_54_fork_io_outputs_1_payload;
    end
    if(inputAll_55_fork_io_outputs_1_ready) begin
      inputAll_55_fork_io_outputs_1_rData <= inputAll_55_fork_io_outputs_1_payload;
    end
    if(inputAll_56_fork_io_outputs_1_ready) begin
      inputAll_56_fork_io_outputs_1_rData <= inputAll_56_fork_io_outputs_1_payload;
    end
    if(inputAll_57_fork_io_outputs_1_ready) begin
      inputAll_57_fork_io_outputs_1_rData <= inputAll_57_fork_io_outputs_1_payload;
    end
    if(inputAll_58_fork_io_outputs_1_ready) begin
      inputAll_58_fork_io_outputs_1_rData <= inputAll_58_fork_io_outputs_1_payload;
    end
    if(inputAll_59_fork_io_outputs_1_ready) begin
      inputAll_59_fork_io_outputs_1_rData <= inputAll_59_fork_io_outputs_1_payload;
    end
    if(inputAll_60_fork_io_outputs_1_ready) begin
      inputAll_60_fork_io_outputs_1_rData <= inputAll_60_fork_io_outputs_1_payload;
    end
    if(inputAll_61_fork_io_outputs_1_ready) begin
      inputAll_61_fork_io_outputs_1_rData <= inputAll_61_fork_io_outputs_1_payload;
    end
    if(inputAll_62_fork_io_outputs_1_ready) begin
      inputAll_62_fork_io_outputs_1_rData <= inputAll_62_fork_io_outputs_1_payload;
    end
    if(inputAll_63_fork_io_outputs_1_ready) begin
      inputAll_63_fork_io_outputs_1_rData <= inputAll_63_fork_io_outputs_1_payload;
    end
    if(inputAll_64_fork_io_outputs_1_ready) begin
      inputAll_64_fork_io_outputs_1_rData <= inputAll_64_fork_io_outputs_1_payload;
    end
    if(inputAll_65_fork_io_outputs_1_ready) begin
      inputAll_65_fork_io_outputs_1_rData <= inputAll_65_fork_io_outputs_1_payload;
    end
    if(inputAll_66_fork_io_outputs_1_ready) begin
      inputAll_66_fork_io_outputs_1_rData <= inputAll_66_fork_io_outputs_1_payload;
    end
    if(inputAll_67_fork_io_outputs_1_ready) begin
      inputAll_67_fork_io_outputs_1_rData <= inputAll_67_fork_io_outputs_1_payload;
    end
    if(inputAll_68_fork_io_outputs_1_ready) begin
      inputAll_68_fork_io_outputs_1_rData <= inputAll_68_fork_io_outputs_1_payload;
    end
    if(inputAll_69_fork_io_outputs_1_ready) begin
      inputAll_69_fork_io_outputs_1_rData <= inputAll_69_fork_io_outputs_1_payload;
    end
    if(inputAll_70_fork_io_outputs_1_ready) begin
      inputAll_70_fork_io_outputs_1_rData <= inputAll_70_fork_io_outputs_1_payload;
    end
    if(inputAll_71_fork_io_outputs_1_ready) begin
      inputAll_71_fork_io_outputs_1_rData <= inputAll_71_fork_io_outputs_1_payload;
    end
    if(inputAll_72_fork_io_outputs_1_ready) begin
      inputAll_72_fork_io_outputs_1_rData <= inputAll_72_fork_io_outputs_1_payload;
    end
    if(inputAll_73_fork_io_outputs_1_ready) begin
      inputAll_73_fork_io_outputs_1_rData <= inputAll_73_fork_io_outputs_1_payload;
    end
    if(inputAll_74_fork_io_outputs_1_ready) begin
      inputAll_74_fork_io_outputs_1_rData <= inputAll_74_fork_io_outputs_1_payload;
    end
    if(inputAll_75_fork_io_outputs_1_ready) begin
      inputAll_75_fork_io_outputs_1_rData <= inputAll_75_fork_io_outputs_1_payload;
    end
    if(inputAll_76_fork_io_outputs_1_ready) begin
      inputAll_76_fork_io_outputs_1_rData <= inputAll_76_fork_io_outputs_1_payload;
    end
    if(inputAll_77_fork_io_outputs_1_ready) begin
      inputAll_77_fork_io_outputs_1_rData <= inputAll_77_fork_io_outputs_1_payload;
    end
    if(inputAll_78_fork_io_outputs_1_ready) begin
      inputAll_78_fork_io_outputs_1_rData <= inputAll_78_fork_io_outputs_1_payload;
    end
    if(inputAll_79_fork_io_outputs_1_ready) begin
      inputAll_79_fork_io_outputs_1_rData <= inputAll_79_fork_io_outputs_1_payload;
    end
    if(inputAll_80_fork_io_outputs_1_ready) begin
      inputAll_80_fork_io_outputs_1_rData <= inputAll_80_fork_io_outputs_1_payload;
    end
    if(inputAll_81_fork_io_outputs_1_ready) begin
      inputAll_81_fork_io_outputs_1_rData <= inputAll_81_fork_io_outputs_1_payload;
    end
    if(inputAll_82_fork_io_outputs_1_ready) begin
      inputAll_82_fork_io_outputs_1_rData <= inputAll_82_fork_io_outputs_1_payload;
    end
    if(inputAll_83_fork_io_outputs_1_ready) begin
      inputAll_83_fork_io_outputs_1_rData <= inputAll_83_fork_io_outputs_1_payload;
    end
    if(inputAll_84_fork_io_outputs_1_ready) begin
      inputAll_84_fork_io_outputs_1_rData <= inputAll_84_fork_io_outputs_1_payload;
    end
    if(inputAll_85_fork_io_outputs_1_ready) begin
      inputAll_85_fork_io_outputs_1_rData <= inputAll_85_fork_io_outputs_1_payload;
    end
    if(inputAll_86_fork_io_outputs_1_ready) begin
      inputAll_86_fork_io_outputs_1_rData <= inputAll_86_fork_io_outputs_1_payload;
    end
    if(inputAll_87_fork_io_outputs_1_ready) begin
      inputAll_87_fork_io_outputs_1_rData <= inputAll_87_fork_io_outputs_1_payload;
    end
    if(inputAll_88_fork_io_outputs_1_ready) begin
      inputAll_88_fork_io_outputs_1_rData <= inputAll_88_fork_io_outputs_1_payload;
    end
    if(inputAll_89_fork_io_outputs_1_ready) begin
      inputAll_89_fork_io_outputs_1_rData <= inputAll_89_fork_io_outputs_1_payload;
    end
    if(inputAll_90_fork_io_outputs_1_ready) begin
      inputAll_90_fork_io_outputs_1_rData <= inputAll_90_fork_io_outputs_1_payload;
    end
    if(inputAll_91_fork_io_outputs_1_ready) begin
      inputAll_91_fork_io_outputs_1_rData <= inputAll_91_fork_io_outputs_1_payload;
    end
    if(inputAll_92_fork_io_outputs_1_ready) begin
      inputAll_92_fork_io_outputs_1_rData <= inputAll_92_fork_io_outputs_1_payload;
    end
    if(inputAll_93_fork_io_outputs_1_ready) begin
      inputAll_93_fork_io_outputs_1_rData <= inputAll_93_fork_io_outputs_1_payload;
    end
    if(inputAll_94_fork_io_outputs_1_ready) begin
      inputAll_94_fork_io_outputs_1_rData <= inputAll_94_fork_io_outputs_1_payload;
    end
    if(inputAll_95_fork_io_outputs_1_ready) begin
      inputAll_95_fork_io_outputs_1_rData <= inputAll_95_fork_io_outputs_1_payload;
    end
    if(inputAll_96_fork_io_outputs_1_ready) begin
      inputAll_96_fork_io_outputs_1_rData <= inputAll_96_fork_io_outputs_1_payload;
    end
    if(inputAll_97_fork_io_outputs_1_ready) begin
      inputAll_97_fork_io_outputs_1_rData <= inputAll_97_fork_io_outputs_1_payload;
    end
    if(inputAll_98_fork_io_outputs_1_ready) begin
      inputAll_98_fork_io_outputs_1_rData <= inputAll_98_fork_io_outputs_1_payload;
    end
    if(inputAll_99_fork_io_outputs_1_ready) begin
      inputAll_99_fork_io_outputs_1_rData <= inputAll_99_fork_io_outputs_1_payload;
    end
    if(inputAll_100_fork_io_outputs_1_ready) begin
      inputAll_100_fork_io_outputs_1_rData <= inputAll_100_fork_io_outputs_1_payload;
    end
    if(inputAll_101_fork_io_outputs_1_ready) begin
      inputAll_101_fork_io_outputs_1_rData <= inputAll_101_fork_io_outputs_1_payload;
    end
    if(inputAll_102_fork_io_outputs_1_ready) begin
      inputAll_102_fork_io_outputs_1_rData <= inputAll_102_fork_io_outputs_1_payload;
    end
    if(inputAll_103_fork_io_outputs_1_ready) begin
      inputAll_103_fork_io_outputs_1_rData <= inputAll_103_fork_io_outputs_1_payload;
    end
    if(inputAll_104_fork_io_outputs_1_ready) begin
      inputAll_104_fork_io_outputs_1_rData <= inputAll_104_fork_io_outputs_1_payload;
    end
    if(inputAll_105_fork_io_outputs_1_ready) begin
      inputAll_105_fork_io_outputs_1_rData <= inputAll_105_fork_io_outputs_1_payload;
    end
    if(inputAll_106_fork_io_outputs_1_ready) begin
      inputAll_106_fork_io_outputs_1_rData <= inputAll_106_fork_io_outputs_1_payload;
    end
    if(inputAll_107_fork_io_outputs_1_ready) begin
      inputAll_107_fork_io_outputs_1_rData <= inputAll_107_fork_io_outputs_1_payload;
    end
    if(inputAll_108_fork_io_outputs_1_ready) begin
      inputAll_108_fork_io_outputs_1_rData <= inputAll_108_fork_io_outputs_1_payload;
    end
    if(inputAll_109_fork_io_outputs_1_ready) begin
      inputAll_109_fork_io_outputs_1_rData <= inputAll_109_fork_io_outputs_1_payload;
    end
    if(inputAll_110_fork_io_outputs_1_ready) begin
      inputAll_110_fork_io_outputs_1_rData <= inputAll_110_fork_io_outputs_1_payload;
    end
    if(inputAll_111_fork_io_outputs_1_ready) begin
      inputAll_111_fork_io_outputs_1_rData <= inputAll_111_fork_io_outputs_1_payload;
    end
    if(inputAll_112_fork_io_outputs_1_ready) begin
      inputAll_112_fork_io_outputs_1_rData <= inputAll_112_fork_io_outputs_1_payload;
    end
    if(inputAll_113_fork_io_outputs_1_ready) begin
      inputAll_113_fork_io_outputs_1_rData <= inputAll_113_fork_io_outputs_1_payload;
    end
    if(inputAll_114_fork_io_outputs_1_ready) begin
      inputAll_114_fork_io_outputs_1_rData <= inputAll_114_fork_io_outputs_1_payload;
    end
    if(inputAll_115_fork_io_outputs_1_ready) begin
      inputAll_115_fork_io_outputs_1_rData <= inputAll_115_fork_io_outputs_1_payload;
    end
    if(inputAll_116_fork_io_outputs_1_ready) begin
      inputAll_116_fork_io_outputs_1_rData <= inputAll_116_fork_io_outputs_1_payload;
    end
    if(inputAll_117_fork_io_outputs_1_ready) begin
      inputAll_117_fork_io_outputs_1_rData <= inputAll_117_fork_io_outputs_1_payload;
    end
    if(inputAll_118_fork_io_outputs_1_ready) begin
      inputAll_118_fork_io_outputs_1_rData <= inputAll_118_fork_io_outputs_1_payload;
    end
    if(inputAll_119_fork_io_outputs_1_ready) begin
      inputAll_119_fork_io_outputs_1_rData <= inputAll_119_fork_io_outputs_1_payload;
    end
    if(inputAll_120_fork_io_outputs_1_ready) begin
      inputAll_120_fork_io_outputs_1_rData <= inputAll_120_fork_io_outputs_1_payload;
    end
    if(inputAll_121_fork_io_outputs_1_ready) begin
      inputAll_121_fork_io_outputs_1_rData <= inputAll_121_fork_io_outputs_1_payload;
    end
    if(inputAll_122_fork_io_outputs_1_ready) begin
      inputAll_122_fork_io_outputs_1_rData <= inputAll_122_fork_io_outputs_1_payload;
    end
    if(inputAll_123_fork_io_outputs_1_ready) begin
      inputAll_123_fork_io_outputs_1_rData <= inputAll_123_fork_io_outputs_1_payload;
    end
    if(inputAll_124_fork_io_outputs_1_ready) begin
      inputAll_124_fork_io_outputs_1_rData <= inputAll_124_fork_io_outputs_1_payload;
    end
    if(inputAll_125_fork_io_outputs_1_ready) begin
      inputAll_125_fork_io_outputs_1_rData <= inputAll_125_fork_io_outputs_1_payload;
    end
    if(inputAll_126_fork_io_outputs_1_ready) begin
      inputAll_126_fork_io_outputs_1_rData <= inputAll_126_fork_io_outputs_1_payload;
    end
    if(inputAll_127_fork_io_outputs_1_ready) begin
      inputAll_127_fork_io_outputs_1_rData <= inputAll_127_fork_io_outputs_1_payload;
    end
  end


endmodule

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

//StreamFork replaced by StreamFork

module StreamFork (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload
);

  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload = io_input_payload;
  assign io_outputs_1_payload = io_input_payload;

endmodule
